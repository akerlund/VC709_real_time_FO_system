library ieee;
use ieee.std_logic_1164.all;
entity chien is
    port(
        a_1     :    in  std_logic_vector(6 downto 0);
        a_2     :    in  std_logic_vector(6 downto 0);
        E     :    out std_logic_vector(126 downto 0)
);
end entity;

architecture arch of chien is
    signal mulr_1_1 : std_logic_vector(6 downto 0);
    signal mulr_2_1 : std_logic_vector(6 downto 0);
    signal mulr_1_2 : std_logic_vector(6 downto 0);
    signal mulr_2_2 : std_logic_vector(6 downto 0);
    signal mulr_1_3 : std_logic_vector(6 downto 0);
    signal mulr_2_3 : std_logic_vector(6 downto 0);
    signal mulr_1_4 : std_logic_vector(6 downto 0);
    signal mulr_2_4 : std_logic_vector(6 downto 0);
    signal mulr_1_5 : std_logic_vector(6 downto 0);
    signal mulr_2_5 : std_logic_vector(6 downto 0);
    signal mulr_1_6 : std_logic_vector(6 downto 0);
    signal mulr_2_6 : std_logic_vector(6 downto 0);
    signal mulr_1_7 : std_logic_vector(6 downto 0);
    signal mulr_2_7 : std_logic_vector(6 downto 0);
    signal mulr_1_8 : std_logic_vector(6 downto 0);
    signal mulr_2_8 : std_logic_vector(6 downto 0);
    signal mulr_1_9 : std_logic_vector(6 downto 0);
    signal mulr_2_9 : std_logic_vector(6 downto 0);
    signal mulr_1_10 : std_logic_vector(6 downto 0);
    signal mulr_2_10 : std_logic_vector(6 downto 0);
    signal mulr_1_11 : std_logic_vector(6 downto 0);
    signal mulr_2_11 : std_logic_vector(6 downto 0);
    signal mulr_1_12 : std_logic_vector(6 downto 0);
    signal mulr_2_12 : std_logic_vector(6 downto 0);
    signal mulr_1_13 : std_logic_vector(6 downto 0);
    signal mulr_2_13 : std_logic_vector(6 downto 0);
    signal mulr_1_14 : std_logic_vector(6 downto 0);
    signal mulr_2_14 : std_logic_vector(6 downto 0);
    signal mulr_1_15 : std_logic_vector(6 downto 0);
    signal mulr_2_15 : std_logic_vector(6 downto 0);
    signal mulr_1_16 : std_logic_vector(6 downto 0);
    signal mulr_2_16 : std_logic_vector(6 downto 0);
    signal mulr_1_17 : std_logic_vector(6 downto 0);
    signal mulr_2_17 : std_logic_vector(6 downto 0);
    signal mulr_1_18 : std_logic_vector(6 downto 0);
    signal mulr_2_18 : std_logic_vector(6 downto 0);
    signal mulr_1_19 : std_logic_vector(6 downto 0);
    signal mulr_2_19 : std_logic_vector(6 downto 0);
    signal mulr_1_20 : std_logic_vector(6 downto 0);
    signal mulr_2_20 : std_logic_vector(6 downto 0);
    signal mulr_1_21 : std_logic_vector(6 downto 0);
    signal mulr_2_21 : std_logic_vector(6 downto 0);
    signal mulr_1_22 : std_logic_vector(6 downto 0);
    signal mulr_2_22 : std_logic_vector(6 downto 0);
    signal mulr_1_23 : std_logic_vector(6 downto 0);
    signal mulr_2_23 : std_logic_vector(6 downto 0);
    signal mulr_1_24 : std_logic_vector(6 downto 0);
    signal mulr_2_24 : std_logic_vector(6 downto 0);
    signal mulr_1_25 : std_logic_vector(6 downto 0);
    signal mulr_2_25 : std_logic_vector(6 downto 0);
    signal mulr_1_26 : std_logic_vector(6 downto 0);
    signal mulr_2_26 : std_logic_vector(6 downto 0);
    signal mulr_1_27 : std_logic_vector(6 downto 0);
    signal mulr_2_27 : std_logic_vector(6 downto 0);
    signal mulr_1_28 : std_logic_vector(6 downto 0);
    signal mulr_2_28 : std_logic_vector(6 downto 0);
    signal mulr_1_29 : std_logic_vector(6 downto 0);
    signal mulr_2_29 : std_logic_vector(6 downto 0);
    signal mulr_1_30 : std_logic_vector(6 downto 0);
    signal mulr_2_30 : std_logic_vector(6 downto 0);
    signal mulr_1_31 : std_logic_vector(6 downto 0);
    signal mulr_2_31 : std_logic_vector(6 downto 0);
    signal mulr_1_32 : std_logic_vector(6 downto 0);
    signal mulr_2_32 : std_logic_vector(6 downto 0);
    signal mulr_1_33 : std_logic_vector(6 downto 0);
    signal mulr_2_33 : std_logic_vector(6 downto 0);
    signal mulr_1_34 : std_logic_vector(6 downto 0);
    signal mulr_2_34 : std_logic_vector(6 downto 0);
    signal mulr_1_35 : std_logic_vector(6 downto 0);
    signal mulr_2_35 : std_logic_vector(6 downto 0);
    signal mulr_1_36 : std_logic_vector(6 downto 0);
    signal mulr_2_36 : std_logic_vector(6 downto 0);
    signal mulr_1_37 : std_logic_vector(6 downto 0);
    signal mulr_2_37 : std_logic_vector(6 downto 0);
    signal mulr_1_38 : std_logic_vector(6 downto 0);
    signal mulr_2_38 : std_logic_vector(6 downto 0);
    signal mulr_1_39 : std_logic_vector(6 downto 0);
    signal mulr_2_39 : std_logic_vector(6 downto 0);
    signal mulr_1_40 : std_logic_vector(6 downto 0);
    signal mulr_2_40 : std_logic_vector(6 downto 0);
    signal mulr_1_41 : std_logic_vector(6 downto 0);
    signal mulr_2_41 : std_logic_vector(6 downto 0);
    signal mulr_1_42 : std_logic_vector(6 downto 0);
    signal mulr_2_42 : std_logic_vector(6 downto 0);
    signal mulr_1_43 : std_logic_vector(6 downto 0);
    signal mulr_2_43 : std_logic_vector(6 downto 0);
    signal mulr_1_44 : std_logic_vector(6 downto 0);
    signal mulr_2_44 : std_logic_vector(6 downto 0);
    signal mulr_1_45 : std_logic_vector(6 downto 0);
    signal mulr_2_45 : std_logic_vector(6 downto 0);
    signal mulr_1_46 : std_logic_vector(6 downto 0);
    signal mulr_2_46 : std_logic_vector(6 downto 0);
    signal mulr_1_47 : std_logic_vector(6 downto 0);
    signal mulr_2_47 : std_logic_vector(6 downto 0);
    signal mulr_1_48 : std_logic_vector(6 downto 0);
    signal mulr_2_48 : std_logic_vector(6 downto 0);
    signal mulr_1_49 : std_logic_vector(6 downto 0);
    signal mulr_2_49 : std_logic_vector(6 downto 0);
    signal mulr_1_50 : std_logic_vector(6 downto 0);
    signal mulr_2_50 : std_logic_vector(6 downto 0);
    signal mulr_1_51 : std_logic_vector(6 downto 0);
    signal mulr_2_51 : std_logic_vector(6 downto 0);
    signal mulr_1_52 : std_logic_vector(6 downto 0);
    signal mulr_2_52 : std_logic_vector(6 downto 0);
    signal mulr_1_53 : std_logic_vector(6 downto 0);
    signal mulr_2_53 : std_logic_vector(6 downto 0);
    signal mulr_1_54 : std_logic_vector(6 downto 0);
    signal mulr_2_54 : std_logic_vector(6 downto 0);
    signal mulr_1_55 : std_logic_vector(6 downto 0);
    signal mulr_2_55 : std_logic_vector(6 downto 0);
    signal mulr_1_56 : std_logic_vector(6 downto 0);
    signal mulr_2_56 : std_logic_vector(6 downto 0);
    signal mulr_1_57 : std_logic_vector(6 downto 0);
    signal mulr_2_57 : std_logic_vector(6 downto 0);
    signal mulr_1_58 : std_logic_vector(6 downto 0);
    signal mulr_2_58 : std_logic_vector(6 downto 0);
    signal mulr_1_59 : std_logic_vector(6 downto 0);
    signal mulr_2_59 : std_logic_vector(6 downto 0);
    signal mulr_1_60 : std_logic_vector(6 downto 0);
    signal mulr_2_60 : std_logic_vector(6 downto 0);
    signal mulr_1_61 : std_logic_vector(6 downto 0);
    signal mulr_2_61 : std_logic_vector(6 downto 0);
    signal mulr_1_62 : std_logic_vector(6 downto 0);
    signal mulr_2_62 : std_logic_vector(6 downto 0);
    signal mulr_1_63 : std_logic_vector(6 downto 0);
    signal mulr_2_63 : std_logic_vector(6 downto 0);
    signal mulr_1_64 : std_logic_vector(6 downto 0);
    signal mulr_2_64 : std_logic_vector(6 downto 0);
    signal mulr_1_65 : std_logic_vector(6 downto 0);
    signal mulr_2_65 : std_logic_vector(6 downto 0);
    signal mulr_1_66 : std_logic_vector(6 downto 0);
    signal mulr_2_66 : std_logic_vector(6 downto 0);
    signal mulr_1_67 : std_logic_vector(6 downto 0);
    signal mulr_2_67 : std_logic_vector(6 downto 0);
    signal mulr_1_68 : std_logic_vector(6 downto 0);
    signal mulr_2_68 : std_logic_vector(6 downto 0);
    signal mulr_1_69 : std_logic_vector(6 downto 0);
    signal mulr_2_69 : std_logic_vector(6 downto 0);
    signal mulr_1_70 : std_logic_vector(6 downto 0);
    signal mulr_2_70 : std_logic_vector(6 downto 0);
    signal mulr_1_71 : std_logic_vector(6 downto 0);
    signal mulr_2_71 : std_logic_vector(6 downto 0);
    signal mulr_1_72 : std_logic_vector(6 downto 0);
    signal mulr_2_72 : std_logic_vector(6 downto 0);
    signal mulr_1_73 : std_logic_vector(6 downto 0);
    signal mulr_2_73 : std_logic_vector(6 downto 0);
    signal mulr_1_74 : std_logic_vector(6 downto 0);
    signal mulr_2_74 : std_logic_vector(6 downto 0);
    signal mulr_1_75 : std_logic_vector(6 downto 0);
    signal mulr_2_75 : std_logic_vector(6 downto 0);
    signal mulr_1_76 : std_logic_vector(6 downto 0);
    signal mulr_2_76 : std_logic_vector(6 downto 0);
    signal mulr_1_77 : std_logic_vector(6 downto 0);
    signal mulr_2_77 : std_logic_vector(6 downto 0);
    signal mulr_1_78 : std_logic_vector(6 downto 0);
    signal mulr_2_78 : std_logic_vector(6 downto 0);
    signal mulr_1_79 : std_logic_vector(6 downto 0);
    signal mulr_2_79 : std_logic_vector(6 downto 0);
    signal mulr_1_80 : std_logic_vector(6 downto 0);
    signal mulr_2_80 : std_logic_vector(6 downto 0);
    signal mulr_1_81 : std_logic_vector(6 downto 0);
    signal mulr_2_81 : std_logic_vector(6 downto 0);
    signal mulr_1_82 : std_logic_vector(6 downto 0);
    signal mulr_2_82 : std_logic_vector(6 downto 0);
    signal mulr_1_83 : std_logic_vector(6 downto 0);
    signal mulr_2_83 : std_logic_vector(6 downto 0);
    signal mulr_1_84 : std_logic_vector(6 downto 0);
    signal mulr_2_84 : std_logic_vector(6 downto 0);
    signal mulr_1_85 : std_logic_vector(6 downto 0);
    signal mulr_2_85 : std_logic_vector(6 downto 0);
    signal mulr_1_86 : std_logic_vector(6 downto 0);
    signal mulr_2_86 : std_logic_vector(6 downto 0);
    signal mulr_1_87 : std_logic_vector(6 downto 0);
    signal mulr_2_87 : std_logic_vector(6 downto 0);
    signal mulr_1_88 : std_logic_vector(6 downto 0);
    signal mulr_2_88 : std_logic_vector(6 downto 0);
    signal mulr_1_89 : std_logic_vector(6 downto 0);
    signal mulr_2_89 : std_logic_vector(6 downto 0);
    signal mulr_1_90 : std_logic_vector(6 downto 0);
    signal mulr_2_90 : std_logic_vector(6 downto 0);
    signal mulr_1_91 : std_logic_vector(6 downto 0);
    signal mulr_2_91 : std_logic_vector(6 downto 0);
    signal mulr_1_92 : std_logic_vector(6 downto 0);
    signal mulr_2_92 : std_logic_vector(6 downto 0);
    signal mulr_1_93 : std_logic_vector(6 downto 0);
    signal mulr_2_93 : std_logic_vector(6 downto 0);
    signal mulr_1_94 : std_logic_vector(6 downto 0);
    signal mulr_2_94 : std_logic_vector(6 downto 0);
    signal mulr_1_95 : std_logic_vector(6 downto 0);
    signal mulr_2_95 : std_logic_vector(6 downto 0);
    signal mulr_1_96 : std_logic_vector(6 downto 0);
    signal mulr_2_96 : std_logic_vector(6 downto 0);
    signal mulr_1_97 : std_logic_vector(6 downto 0);
    signal mulr_2_97 : std_logic_vector(6 downto 0);
    signal mulr_1_98 : std_logic_vector(6 downto 0);
    signal mulr_2_98 : std_logic_vector(6 downto 0);
    signal mulr_1_99 : std_logic_vector(6 downto 0);
    signal mulr_2_99 : std_logic_vector(6 downto 0);
    signal mulr_1_100 : std_logic_vector(6 downto 0);
    signal mulr_2_100 : std_logic_vector(6 downto 0);
    signal mulr_1_101 : std_logic_vector(6 downto 0);
    signal mulr_2_101 : std_logic_vector(6 downto 0);
    signal mulr_1_102 : std_logic_vector(6 downto 0);
    signal mulr_2_102 : std_logic_vector(6 downto 0);
    signal mulr_1_103 : std_logic_vector(6 downto 0);
    signal mulr_2_103 : std_logic_vector(6 downto 0);
    signal mulr_1_104 : std_logic_vector(6 downto 0);
    signal mulr_2_104 : std_logic_vector(6 downto 0);
    signal mulr_1_105 : std_logic_vector(6 downto 0);
    signal mulr_2_105 : std_logic_vector(6 downto 0);
    signal mulr_1_106 : std_logic_vector(6 downto 0);
    signal mulr_2_106 : std_logic_vector(6 downto 0);
    signal mulr_1_107 : std_logic_vector(6 downto 0);
    signal mulr_2_107 : std_logic_vector(6 downto 0);
    signal mulr_1_108 : std_logic_vector(6 downto 0);
    signal mulr_2_108 : std_logic_vector(6 downto 0);
    signal mulr_1_109 : std_logic_vector(6 downto 0);
    signal mulr_2_109 : std_logic_vector(6 downto 0);
    signal mulr_1_110 : std_logic_vector(6 downto 0);
    signal mulr_2_110 : std_logic_vector(6 downto 0);
    signal mulr_1_111 : std_logic_vector(6 downto 0);
    signal mulr_2_111 : std_logic_vector(6 downto 0);
    signal mulr_1_112 : std_logic_vector(6 downto 0);
    signal mulr_2_112 : std_logic_vector(6 downto 0);
    signal mulr_1_113 : std_logic_vector(6 downto 0);
    signal mulr_2_113 : std_logic_vector(6 downto 0);
    signal mulr_1_114 : std_logic_vector(6 downto 0);
    signal mulr_2_114 : std_logic_vector(6 downto 0);
    signal mulr_1_115 : std_logic_vector(6 downto 0);
    signal mulr_2_115 : std_logic_vector(6 downto 0);
    signal mulr_1_116 : std_logic_vector(6 downto 0);
    signal mulr_2_116 : std_logic_vector(6 downto 0);
    signal mulr_1_117 : std_logic_vector(6 downto 0);
    signal mulr_2_117 : std_logic_vector(6 downto 0);
    signal mulr_1_118 : std_logic_vector(6 downto 0);
    signal mulr_2_118 : std_logic_vector(6 downto 0);
    signal mulr_1_119 : std_logic_vector(6 downto 0);
    signal mulr_2_119 : std_logic_vector(6 downto 0);
    signal mulr_1_120 : std_logic_vector(6 downto 0);
    signal mulr_2_120 : std_logic_vector(6 downto 0);
    signal mulr_1_121 : std_logic_vector(6 downto 0);
    signal mulr_2_121 : std_logic_vector(6 downto 0);
    signal mulr_1_122 : std_logic_vector(6 downto 0);
    signal mulr_2_122 : std_logic_vector(6 downto 0);
    signal mulr_1_123 : std_logic_vector(6 downto 0);
    signal mulr_2_123 : std_logic_vector(6 downto 0);
    signal mulr_1_124 : std_logic_vector(6 downto 0);
    signal mulr_2_124 : std_logic_vector(6 downto 0);
    signal mulr_1_125 : std_logic_vector(6 downto 0);
    signal mulr_2_125 : std_logic_vector(6 downto 0);
    signal mulr_1_126 : std_logic_vector(6 downto 0);
    signal mulr_2_126 : std_logic_vector(6 downto 0);
    signal mulr_1_127 : std_logic_vector(6 downto 0);
    signal mulr_2_127 : std_logic_vector(6 downto 0);
    signal sumr_1 : std_logic_vector(6 downto 0);
    signal sumr_2 : std_logic_vector(6 downto 0);
    signal sumr_3 : std_logic_vector(6 downto 0);
    signal sumr_4 : std_logic_vector(6 downto 0);
    signal sumr_5 : std_logic_vector(6 downto 0);
    signal sumr_6 : std_logic_vector(6 downto 0);
    signal sumr_7 : std_logic_vector(6 downto 0);
    signal sumr_8 : std_logic_vector(6 downto 0);
    signal sumr_9 : std_logic_vector(6 downto 0);
    signal sumr_10 : std_logic_vector(6 downto 0);
    signal sumr_11 : std_logic_vector(6 downto 0);
    signal sumr_12 : std_logic_vector(6 downto 0);
    signal sumr_13 : std_logic_vector(6 downto 0);
    signal sumr_14 : std_logic_vector(6 downto 0);
    signal sumr_15 : std_logic_vector(6 downto 0);
    signal sumr_16 : std_logic_vector(6 downto 0);
    signal sumr_17 : std_logic_vector(6 downto 0);
    signal sumr_18 : std_logic_vector(6 downto 0);
    signal sumr_19 : std_logic_vector(6 downto 0);
    signal sumr_20 : std_logic_vector(6 downto 0);
    signal sumr_21 : std_logic_vector(6 downto 0);
    signal sumr_22 : std_logic_vector(6 downto 0);
    signal sumr_23 : std_logic_vector(6 downto 0);
    signal sumr_24 : std_logic_vector(6 downto 0);
    signal sumr_25 : std_logic_vector(6 downto 0);
    signal sumr_26 : std_logic_vector(6 downto 0);
    signal sumr_27 : std_logic_vector(6 downto 0);
    signal sumr_28 : std_logic_vector(6 downto 0);
    signal sumr_29 : std_logic_vector(6 downto 0);
    signal sumr_30 : std_logic_vector(6 downto 0);
    signal sumr_31 : std_logic_vector(6 downto 0);
    signal sumr_32 : std_logic_vector(6 downto 0);
    signal sumr_33 : std_logic_vector(6 downto 0);
    signal sumr_34 : std_logic_vector(6 downto 0);
    signal sumr_35 : std_logic_vector(6 downto 0);
    signal sumr_36 : std_logic_vector(6 downto 0);
    signal sumr_37 : std_logic_vector(6 downto 0);
    signal sumr_38 : std_logic_vector(6 downto 0);
    signal sumr_39 : std_logic_vector(6 downto 0);
    signal sumr_40 : std_logic_vector(6 downto 0);
    signal sumr_41 : std_logic_vector(6 downto 0);
    signal sumr_42 : std_logic_vector(6 downto 0);
    signal sumr_43 : std_logic_vector(6 downto 0);
    signal sumr_44 : std_logic_vector(6 downto 0);
    signal sumr_45 : std_logic_vector(6 downto 0);
    signal sumr_46 : std_logic_vector(6 downto 0);
    signal sumr_47 : std_logic_vector(6 downto 0);
    signal sumr_48 : std_logic_vector(6 downto 0);
    signal sumr_49 : std_logic_vector(6 downto 0);
    signal sumr_50 : std_logic_vector(6 downto 0);
    signal sumr_51 : std_logic_vector(6 downto 0);
    signal sumr_52 : std_logic_vector(6 downto 0);
    signal sumr_53 : std_logic_vector(6 downto 0);
    signal sumr_54 : std_logic_vector(6 downto 0);
    signal sumr_55 : std_logic_vector(6 downto 0);
    signal sumr_56 : std_logic_vector(6 downto 0);
    signal sumr_57 : std_logic_vector(6 downto 0);
    signal sumr_58 : std_logic_vector(6 downto 0);
    signal sumr_59 : std_logic_vector(6 downto 0);
    signal sumr_60 : std_logic_vector(6 downto 0);
    signal sumr_61 : std_logic_vector(6 downto 0);
    signal sumr_62 : std_logic_vector(6 downto 0);
    signal sumr_63 : std_logic_vector(6 downto 0);
    signal sumr_64 : std_logic_vector(6 downto 0);
    signal sumr_65 : std_logic_vector(6 downto 0);
    signal sumr_66 : std_logic_vector(6 downto 0);
    signal sumr_67 : std_logic_vector(6 downto 0);
    signal sumr_68 : std_logic_vector(6 downto 0);
    signal sumr_69 : std_logic_vector(6 downto 0);
    signal sumr_70 : std_logic_vector(6 downto 0);
    signal sumr_71 : std_logic_vector(6 downto 0);
    signal sumr_72 : std_logic_vector(6 downto 0);
    signal sumr_73 : std_logic_vector(6 downto 0);
    signal sumr_74 : std_logic_vector(6 downto 0);
    signal sumr_75 : std_logic_vector(6 downto 0);
    signal sumr_76 : std_logic_vector(6 downto 0);
    signal sumr_77 : std_logic_vector(6 downto 0);
    signal sumr_78 : std_logic_vector(6 downto 0);
    signal sumr_79 : std_logic_vector(6 downto 0);
    signal sumr_80 : std_logic_vector(6 downto 0);
    signal sumr_81 : std_logic_vector(6 downto 0);
    signal sumr_82 : std_logic_vector(6 downto 0);
    signal sumr_83 : std_logic_vector(6 downto 0);
    signal sumr_84 : std_logic_vector(6 downto 0);
    signal sumr_85 : std_logic_vector(6 downto 0);
    signal sumr_86 : std_logic_vector(6 downto 0);
    signal sumr_87 : std_logic_vector(6 downto 0);
    signal sumr_88 : std_logic_vector(6 downto 0);
    signal sumr_89 : std_logic_vector(6 downto 0);
    signal sumr_90 : std_logic_vector(6 downto 0);
    signal sumr_91 : std_logic_vector(6 downto 0);
    signal sumr_92 : std_logic_vector(6 downto 0);
    signal sumr_93 : std_logic_vector(6 downto 0);
    signal sumr_94 : std_logic_vector(6 downto 0);
    signal sumr_95 : std_logic_vector(6 downto 0);
    signal sumr_96 : std_logic_vector(6 downto 0);
    signal sumr_97 : std_logic_vector(6 downto 0);
    signal sumr_98 : std_logic_vector(6 downto 0);
    signal sumr_99 : std_logic_vector(6 downto 0);
    signal sumr_100 : std_logic_vector(6 downto 0);
    signal sumr_101 : std_logic_vector(6 downto 0);
    signal sumr_102 : std_logic_vector(6 downto 0);
    signal sumr_103 : std_logic_vector(6 downto 0);
    signal sumr_104 : std_logic_vector(6 downto 0);
    signal sumr_105 : std_logic_vector(6 downto 0);
    signal sumr_106 : std_logic_vector(6 downto 0);
    signal sumr_107 : std_logic_vector(6 downto 0);
    signal sumr_108 : std_logic_vector(6 downto 0);
    signal sumr_109 : std_logic_vector(6 downto 0);
    signal sumr_110 : std_logic_vector(6 downto 0);
    signal sumr_111 : std_logic_vector(6 downto 0);
    signal sumr_112 : std_logic_vector(6 downto 0);
    signal sumr_113 : std_logic_vector(6 downto 0);
    signal sumr_114 : std_logic_vector(6 downto 0);
    signal sumr_115 : std_logic_vector(6 downto 0);
    signal sumr_116 : std_logic_vector(6 downto 0);
    signal sumr_117 : std_logic_vector(6 downto 0);
    signal sumr_118 : std_logic_vector(6 downto 0);
    signal sumr_119 : std_logic_vector(6 downto 0);
    signal sumr_120 : std_logic_vector(6 downto 0);
    signal sumr_121 : std_logic_vector(6 downto 0);
    signal sumr_122 : std_logic_vector(6 downto 0);
    signal sumr_123 : std_logic_vector(6 downto 0);
    signal sumr_124 : std_logic_vector(6 downto 0);
    signal sumr_125 : std_logic_vector(6 downto 0);
    signal sumr_126 : std_logic_vector(6 downto 0);
    signal sumr_127 : std_logic_vector(6 downto 0);
begin

mulr_1_1<=a_1;
mulc_2_1 : entity work.gfmul
port map(
a=>a_2,
b=>"0000010",
X=>mulr_2_1);

mulr_1_2<=a_1;
mulc_2_2 : entity work.gfmul
port map(
a=>a_2,
b=>"0000100",
X=>mulr_2_2);

mulr_1_3<=a_1;
mulc_2_3 : entity work.gfmul
port map(
a=>a_2,
b=>"0001000",
X=>mulr_2_3);

mulr_1_4<=a_1;
mulc_2_4 : entity work.gfmul
port map(
a=>a_2,
b=>"0010000",
X=>mulr_2_4);

mulr_1_5<=a_1;
mulc_2_5 : entity work.gfmul
port map(
a=>a_2,
b=>"0100000",
X=>mulr_2_5);

mulr_1_6<=a_1;
mulc_2_6 : entity work.gfmul
port map(
a=>a_2,
b=>"1000000",
X=>mulr_2_6);

mulr_1_7<=a_1;
mulc_2_7 : entity work.gfmul
port map(
a=>a_2,
b=>"0001001",
X=>mulr_2_7);

mulr_1_8<=a_1;
mulc_2_8 : entity work.gfmul
port map(
a=>a_2,
b=>"0010010",
X=>mulr_2_8);

mulr_1_9<=a_1;
mulc_2_9 : entity work.gfmul
port map(
a=>a_2,
b=>"0100100",
X=>mulr_2_9);

mulr_1_10<=a_1;
mulc_2_10 : entity work.gfmul
port map(
a=>a_2,
b=>"1001000",
X=>mulr_2_10);

mulr_1_11<=a_1;
mulc_2_11 : entity work.gfmul
port map(
a=>a_2,
b=>"0011001",
X=>mulr_2_11);

mulr_1_12<=a_1;
mulc_2_12 : entity work.gfmul
port map(
a=>a_2,
b=>"0110010",
X=>mulr_2_12);

mulr_1_13<=a_1;
mulc_2_13 : entity work.gfmul
port map(
a=>a_2,
b=>"1100100",
X=>mulr_2_13);

mulr_1_14<=a_1;
mulc_2_14 : entity work.gfmul
port map(
a=>a_2,
b=>"1000001",
X=>mulr_2_14);

mulr_1_15<=a_1;
mulc_2_15 : entity work.gfmul
port map(
a=>a_2,
b=>"0001011",
X=>mulr_2_15);

mulr_1_16<=a_1;
mulc_2_16 : entity work.gfmul
port map(
a=>a_2,
b=>"0010110",
X=>mulr_2_16);

mulr_1_17<=a_1;
mulc_2_17 : entity work.gfmul
port map(
a=>a_2,
b=>"0101100",
X=>mulr_2_17);

mulr_1_18<=a_1;
mulc_2_18 : entity work.gfmul
port map(
a=>a_2,
b=>"1011000",
X=>mulr_2_18);

mulr_1_19<=a_1;
mulc_2_19 : entity work.gfmul
port map(
a=>a_2,
b=>"0111001",
X=>mulr_2_19);

mulr_1_20<=a_1;
mulc_2_20 : entity work.gfmul
port map(
a=>a_2,
b=>"1110010",
X=>mulr_2_20);

mulr_1_21<=a_1;
mulc_2_21 : entity work.gfmul
port map(
a=>a_2,
b=>"1101101",
X=>mulr_2_21);

mulr_1_22<=a_1;
mulc_2_22 : entity work.gfmul
port map(
a=>a_2,
b=>"1010011",
X=>mulr_2_22);

mulr_1_23<=a_1;
mulc_2_23 : entity work.gfmul
port map(
a=>a_2,
b=>"0101111",
X=>mulr_2_23);

mulr_1_24<=a_1;
mulc_2_24 : entity work.gfmul
port map(
a=>a_2,
b=>"1011110",
X=>mulr_2_24);

mulr_1_25<=a_1;
mulc_2_25 : entity work.gfmul
port map(
a=>a_2,
b=>"0110101",
X=>mulr_2_25);

mulr_1_26<=a_1;
mulc_2_26 : entity work.gfmul
port map(
a=>a_2,
b=>"1101010",
X=>mulr_2_26);

mulr_1_27<=a_1;
mulc_2_27 : entity work.gfmul
port map(
a=>a_2,
b=>"1011101",
X=>mulr_2_27);

mulr_1_28<=a_1;
mulc_2_28 : entity work.gfmul
port map(
a=>a_2,
b=>"0110011",
X=>mulr_2_28);

mulr_1_29<=a_1;
mulc_2_29 : entity work.gfmul
port map(
a=>a_2,
b=>"1100110",
X=>mulr_2_29);

mulr_1_30<=a_1;
mulc_2_30 : entity work.gfmul
port map(
a=>a_2,
b=>"1000101",
X=>mulr_2_30);

mulr_1_31<=a_1;
mulc_2_31 : entity work.gfmul
port map(
a=>a_2,
b=>"0000011",
X=>mulr_2_31);

mulr_1_32<=a_1;
mulc_2_32 : entity work.gfmul
port map(
a=>a_2,
b=>"0000110",
X=>mulr_2_32);

mulr_1_33<=a_1;
mulc_2_33 : entity work.gfmul
port map(
a=>a_2,
b=>"0001100",
X=>mulr_2_33);

mulr_1_34<=a_1;
mulc_2_34 : entity work.gfmul
port map(
a=>a_2,
b=>"0011000",
X=>mulr_2_34);

mulr_1_35<=a_1;
mulc_2_35 : entity work.gfmul
port map(
a=>a_2,
b=>"0110000",
X=>mulr_2_35);

mulr_1_36<=a_1;
mulc_2_36 : entity work.gfmul
port map(
a=>a_2,
b=>"1100000",
X=>mulr_2_36);

mulr_1_37<=a_1;
mulc_2_37 : entity work.gfmul
port map(
a=>a_2,
b=>"1001001",
X=>mulr_2_37);

mulr_1_38<=a_1;
mulc_2_38 : entity work.gfmul
port map(
a=>a_2,
b=>"0011011",
X=>mulr_2_38);

mulr_1_39<=a_1;
mulc_2_39 : entity work.gfmul
port map(
a=>a_2,
b=>"0110110",
X=>mulr_2_39);

mulr_1_40<=a_1;
mulc_2_40 : entity work.gfmul
port map(
a=>a_2,
b=>"1101100",
X=>mulr_2_40);

mulr_1_41<=a_1;
mulc_2_41 : entity work.gfmul
port map(
a=>a_2,
b=>"1010001",
X=>mulr_2_41);

mulr_1_42<=a_1;
mulc_2_42 : entity work.gfmul
port map(
a=>a_2,
b=>"0101011",
X=>mulr_2_42);

mulr_1_43<=a_1;
mulc_2_43 : entity work.gfmul
port map(
a=>a_2,
b=>"1010110",
X=>mulr_2_43);

mulr_1_44<=a_1;
mulc_2_44 : entity work.gfmul
port map(
a=>a_2,
b=>"0100101",
X=>mulr_2_44);

mulr_1_45<=a_1;
mulc_2_45 : entity work.gfmul
port map(
a=>a_2,
b=>"1001010",
X=>mulr_2_45);

mulr_1_46<=a_1;
mulc_2_46 : entity work.gfmul
port map(
a=>a_2,
b=>"0011101",
X=>mulr_2_46);

mulr_1_47<=a_1;
mulc_2_47 : entity work.gfmul
port map(
a=>a_2,
b=>"0111010",
X=>mulr_2_47);

mulr_1_48<=a_1;
mulc_2_48 : entity work.gfmul
port map(
a=>a_2,
b=>"1110100",
X=>mulr_2_48);

mulr_1_49<=a_1;
mulc_2_49 : entity work.gfmul
port map(
a=>a_2,
b=>"1100001",
X=>mulr_2_49);

mulr_1_50<=a_1;
mulc_2_50 : entity work.gfmul
port map(
a=>a_2,
b=>"1001011",
X=>mulr_2_50);

mulr_1_51<=a_1;
mulc_2_51 : entity work.gfmul
port map(
a=>a_2,
b=>"0011111",
X=>mulr_2_51);

mulr_1_52<=a_1;
mulc_2_52 : entity work.gfmul
port map(
a=>a_2,
b=>"0111110",
X=>mulr_2_52);

mulr_1_53<=a_1;
mulc_2_53 : entity work.gfmul
port map(
a=>a_2,
b=>"1111100",
X=>mulr_2_53);

mulr_1_54<=a_1;
mulc_2_54 : entity work.gfmul
port map(
a=>a_2,
b=>"1110001",
X=>mulr_2_54);

mulr_1_55<=a_1;
mulc_2_55 : entity work.gfmul
port map(
a=>a_2,
b=>"1101011",
X=>mulr_2_55);

mulr_1_56<=a_1;
mulc_2_56 : entity work.gfmul
port map(
a=>a_2,
b=>"1011111",
X=>mulr_2_56);

mulr_1_57<=a_1;
mulc_2_57 : entity work.gfmul
port map(
a=>a_2,
b=>"0110111",
X=>mulr_2_57);

mulr_1_58<=a_1;
mulc_2_58 : entity work.gfmul
port map(
a=>a_2,
b=>"1101110",
X=>mulr_2_58);

mulr_1_59<=a_1;
mulc_2_59 : entity work.gfmul
port map(
a=>a_2,
b=>"1010101",
X=>mulr_2_59);

mulr_1_60<=a_1;
mulc_2_60 : entity work.gfmul
port map(
a=>a_2,
b=>"0100011",
X=>mulr_2_60);

mulr_1_61<=a_1;
mulc_2_61 : entity work.gfmul
port map(
a=>a_2,
b=>"1000110",
X=>mulr_2_61);

mulr_1_62<=a_1;
mulc_2_62 : entity work.gfmul
port map(
a=>a_2,
b=>"0000101",
X=>mulr_2_62);

mulr_1_63<=a_1;
mulc_2_63 : entity work.gfmul
port map(
a=>a_2,
b=>"0001010",
X=>mulr_2_63);

mulr_1_64<=a_1;
mulc_2_64 : entity work.gfmul
port map(
a=>a_2,
b=>"0010100",
X=>mulr_2_64);

mulr_1_65<=a_1;
mulc_2_65 : entity work.gfmul
port map(
a=>a_2,
b=>"0101000",
X=>mulr_2_65);

mulr_1_66<=a_1;
mulc_2_66 : entity work.gfmul
port map(
a=>a_2,
b=>"1010000",
X=>mulr_2_66);

mulr_1_67<=a_1;
mulc_2_67 : entity work.gfmul
port map(
a=>a_2,
b=>"0101001",
X=>mulr_2_67);

mulr_1_68<=a_1;
mulc_2_68 : entity work.gfmul
port map(
a=>a_2,
b=>"1010010",
X=>mulr_2_68);

mulr_1_69<=a_1;
mulc_2_69 : entity work.gfmul
port map(
a=>a_2,
b=>"0101101",
X=>mulr_2_69);

mulr_1_70<=a_1;
mulc_2_70 : entity work.gfmul
port map(
a=>a_2,
b=>"1011010",
X=>mulr_2_70);

mulr_1_71<=a_1;
mulc_2_71 : entity work.gfmul
port map(
a=>a_2,
b=>"0111101",
X=>mulr_2_71);

mulr_1_72<=a_1;
mulc_2_72 : entity work.gfmul
port map(
a=>a_2,
b=>"1111010",
X=>mulr_2_72);

mulr_1_73<=a_1;
mulc_2_73 : entity work.gfmul
port map(
a=>a_2,
b=>"1111101",
X=>mulr_2_73);

mulr_1_74<=a_1;
mulc_2_74 : entity work.gfmul
port map(
a=>a_2,
b=>"1110011",
X=>mulr_2_74);

mulr_1_75<=a_1;
mulc_2_75 : entity work.gfmul
port map(
a=>a_2,
b=>"1101111",
X=>mulr_2_75);

mulr_1_76<=a_1;
mulc_2_76 : entity work.gfmul
port map(
a=>a_2,
b=>"1010111",
X=>mulr_2_76);

mulr_1_77<=a_1;
mulc_2_77 : entity work.gfmul
port map(
a=>a_2,
b=>"0100111",
X=>mulr_2_77);

mulr_1_78<=a_1;
mulc_2_78 : entity work.gfmul
port map(
a=>a_2,
b=>"1001110",
X=>mulr_2_78);

mulr_1_79<=a_1;
mulc_2_79 : entity work.gfmul
port map(
a=>a_2,
b=>"0010101",
X=>mulr_2_79);

mulr_1_80<=a_1;
mulc_2_80 : entity work.gfmul
port map(
a=>a_2,
b=>"0101010",
X=>mulr_2_80);

mulr_1_81<=a_1;
mulc_2_81 : entity work.gfmul
port map(
a=>a_2,
b=>"1010100",
X=>mulr_2_81);

mulr_1_82<=a_1;
mulc_2_82 : entity work.gfmul
port map(
a=>a_2,
b=>"0100001",
X=>mulr_2_82);

mulr_1_83<=a_1;
mulc_2_83 : entity work.gfmul
port map(
a=>a_2,
b=>"1000010",
X=>mulr_2_83);

mulr_1_84<=a_1;
mulc_2_84 : entity work.gfmul
port map(
a=>a_2,
b=>"0001101",
X=>mulr_2_84);

mulr_1_85<=a_1;
mulc_2_85 : entity work.gfmul
port map(
a=>a_2,
b=>"0011010",
X=>mulr_2_85);

mulr_1_86<=a_1;
mulc_2_86 : entity work.gfmul
port map(
a=>a_2,
b=>"0110100",
X=>mulr_2_86);

mulr_1_87<=a_1;
mulc_2_87 : entity work.gfmul
port map(
a=>a_2,
b=>"1101000",
X=>mulr_2_87);

mulr_1_88<=a_1;
mulc_2_88 : entity work.gfmul
port map(
a=>a_2,
b=>"1011001",
X=>mulr_2_88);

mulr_1_89<=a_1;
mulc_2_89 : entity work.gfmul
port map(
a=>a_2,
b=>"0111011",
X=>mulr_2_89);

mulr_1_90<=a_1;
mulc_2_90 : entity work.gfmul
port map(
a=>a_2,
b=>"1110110",
X=>mulr_2_90);

mulr_1_91<=a_1;
mulc_2_91 : entity work.gfmul
port map(
a=>a_2,
b=>"1100101",
X=>mulr_2_91);

mulr_1_92<=a_1;
mulc_2_92 : entity work.gfmul
port map(
a=>a_2,
b=>"1000011",
X=>mulr_2_92);

mulr_1_93<=a_1;
mulc_2_93 : entity work.gfmul
port map(
a=>a_2,
b=>"0001111",
X=>mulr_2_93);

mulr_1_94<=a_1;
mulc_2_94 : entity work.gfmul
port map(
a=>a_2,
b=>"0011110",
X=>mulr_2_94);

mulr_1_95<=a_1;
mulc_2_95 : entity work.gfmul
port map(
a=>a_2,
b=>"0111100",
X=>mulr_2_95);

mulr_1_96<=a_1;
mulc_2_96 : entity work.gfmul
port map(
a=>a_2,
b=>"1111000",
X=>mulr_2_96);

mulr_1_97<=a_1;
mulc_2_97 : entity work.gfmul
port map(
a=>a_2,
b=>"1111001",
X=>mulr_2_97);

mulr_1_98<=a_1;
mulc_2_98 : entity work.gfmul
port map(
a=>a_2,
b=>"1111011",
X=>mulr_2_98);

mulr_1_99<=a_1;
mulc_2_99 : entity work.gfmul
port map(
a=>a_2,
b=>"1111111",
X=>mulr_2_99);

mulr_1_100<=a_1;
mulc_2_100 : entity work.gfmul
port map(
a=>a_2,
b=>"1110111",
X=>mulr_2_100);

mulr_1_101<=a_1;
mulc_2_101 : entity work.gfmul
port map(
a=>a_2,
b=>"1100111",
X=>mulr_2_101);

mulr_1_102<=a_1;
mulc_2_102 : entity work.gfmul
port map(
a=>a_2,
b=>"1000111",
X=>mulr_2_102);

mulr_1_103<=a_1;
mulc_2_103 : entity work.gfmul
port map(
a=>a_2,
b=>"0000111",
X=>mulr_2_103);

mulr_1_104<=a_1;
mulc_2_104 : entity work.gfmul
port map(
a=>a_2,
b=>"0001110",
X=>mulr_2_104);

mulr_1_105<=a_1;
mulc_2_105 : entity work.gfmul
port map(
a=>a_2,
b=>"0011100",
X=>mulr_2_105);

mulr_1_106<=a_1;
mulc_2_106 : entity work.gfmul
port map(
a=>a_2,
b=>"0111000",
X=>mulr_2_106);

mulr_1_107<=a_1;
mulc_2_107 : entity work.gfmul
port map(
a=>a_2,
b=>"1110000",
X=>mulr_2_107);

mulr_1_108<=a_1;
mulc_2_108 : entity work.gfmul
port map(
a=>a_2,
b=>"1101001",
X=>mulr_2_108);

mulr_1_109<=a_1;
mulc_2_109 : entity work.gfmul
port map(
a=>a_2,
b=>"1011011",
X=>mulr_2_109);

mulr_1_110<=a_1;
mulc_2_110 : entity work.gfmul
port map(
a=>a_2,
b=>"0111111",
X=>mulr_2_110);

mulr_1_111<=a_1;
mulc_2_111 : entity work.gfmul
port map(
a=>a_2,
b=>"1111110",
X=>mulr_2_111);

mulr_1_112<=a_1;
mulc_2_112 : entity work.gfmul
port map(
a=>a_2,
b=>"1110101",
X=>mulr_2_112);

mulr_1_113<=a_1;
mulc_2_113 : entity work.gfmul
port map(
a=>a_2,
b=>"1100011",
X=>mulr_2_113);

mulr_1_114<=a_1;
mulc_2_114 : entity work.gfmul
port map(
a=>a_2,
b=>"1001111",
X=>mulr_2_114);

mulr_1_115<=a_1;
mulc_2_115 : entity work.gfmul
port map(
a=>a_2,
b=>"0010111",
X=>mulr_2_115);

mulr_1_116<=a_1;
mulc_2_116 : entity work.gfmul
port map(
a=>a_2,
b=>"0101110",
X=>mulr_2_116);

mulr_1_117<=a_1;
mulc_2_117 : entity work.gfmul
port map(
a=>a_2,
b=>"1011100",
X=>mulr_2_117);

mulr_1_118<=a_1;
mulc_2_118 : entity work.gfmul
port map(
a=>a_2,
b=>"0110001",
X=>mulr_2_118);

mulr_1_119<=a_1;
mulc_2_119 : entity work.gfmul
port map(
a=>a_2,
b=>"1100010",
X=>mulr_2_119);

mulr_1_120<=a_1;
mulc_2_120 : entity work.gfmul
port map(
a=>a_2,
b=>"1001101",
X=>mulr_2_120);

mulr_1_121<=a_1;
mulc_2_121 : entity work.gfmul
port map(
a=>a_2,
b=>"0010011",
X=>mulr_2_121);

mulr_1_122<=a_1;
mulc_2_122 : entity work.gfmul
port map(
a=>a_2,
b=>"0100110",
X=>mulr_2_122);

mulr_1_123<=a_1;
mulc_2_123 : entity work.gfmul
port map(
a=>a_2,
b=>"1001100",
X=>mulr_2_123);

mulr_1_124<=a_1;
mulc_2_124 : entity work.gfmul
port map(
a=>a_2,
b=>"0010001",
X=>mulr_2_124);

mulr_1_125<=a_1;
mulc_2_125 : entity work.gfmul
port map(
a=>a_2,
b=>"0100010",
X=>mulr_2_125);

mulr_1_126<=a_1;
mulc_2_126 : entity work.gfmul
port map(
a=>a_2,
b=>"1000100",
X=>mulr_2_126);

mulr_1_127<=a_1;
mulc_2_127 : entity work.gfmul
port map(
a=>a_2,
b=>"0000001",
X=>mulr_2_127);

sumr_1<= mulr_1_1 xor mulr_2_1;
sumr_2<= mulr_1_2 xor mulr_2_2;
sumr_3<= mulr_1_3 xor mulr_2_3;
sumr_4<= mulr_1_4 xor mulr_2_4;
sumr_5<= mulr_1_5 xor mulr_2_5;
sumr_6<= mulr_1_6 xor mulr_2_6;
sumr_7<= mulr_1_7 xor mulr_2_7;
sumr_8<= mulr_1_8 xor mulr_2_8;
sumr_9<= mulr_1_9 xor mulr_2_9;
sumr_10<= mulr_1_10 xor mulr_2_10;
sumr_11<= mulr_1_11 xor mulr_2_11;
sumr_12<= mulr_1_12 xor mulr_2_12;
sumr_13<= mulr_1_13 xor mulr_2_13;
sumr_14<= mulr_1_14 xor mulr_2_14;
sumr_15<= mulr_1_15 xor mulr_2_15;
sumr_16<= mulr_1_16 xor mulr_2_16;
sumr_17<= mulr_1_17 xor mulr_2_17;
sumr_18<= mulr_1_18 xor mulr_2_18;
sumr_19<= mulr_1_19 xor mulr_2_19;
sumr_20<= mulr_1_20 xor mulr_2_20;
sumr_21<= mulr_1_21 xor mulr_2_21;
sumr_22<= mulr_1_22 xor mulr_2_22;
sumr_23<= mulr_1_23 xor mulr_2_23;
sumr_24<= mulr_1_24 xor mulr_2_24;
sumr_25<= mulr_1_25 xor mulr_2_25;
sumr_26<= mulr_1_26 xor mulr_2_26;
sumr_27<= mulr_1_27 xor mulr_2_27;
sumr_28<= mulr_1_28 xor mulr_2_28;
sumr_29<= mulr_1_29 xor mulr_2_29;
sumr_30<= mulr_1_30 xor mulr_2_30;
sumr_31<= mulr_1_31 xor mulr_2_31;
sumr_32<= mulr_1_32 xor mulr_2_32;
sumr_33<= mulr_1_33 xor mulr_2_33;
sumr_34<= mulr_1_34 xor mulr_2_34;
sumr_35<= mulr_1_35 xor mulr_2_35;
sumr_36<= mulr_1_36 xor mulr_2_36;
sumr_37<= mulr_1_37 xor mulr_2_37;
sumr_38<= mulr_1_38 xor mulr_2_38;
sumr_39<= mulr_1_39 xor mulr_2_39;
sumr_40<= mulr_1_40 xor mulr_2_40;
sumr_41<= mulr_1_41 xor mulr_2_41;
sumr_42<= mulr_1_42 xor mulr_2_42;
sumr_43<= mulr_1_43 xor mulr_2_43;
sumr_44<= mulr_1_44 xor mulr_2_44;
sumr_45<= mulr_1_45 xor mulr_2_45;
sumr_46<= mulr_1_46 xor mulr_2_46;
sumr_47<= mulr_1_47 xor mulr_2_47;
sumr_48<= mulr_1_48 xor mulr_2_48;
sumr_49<= mulr_1_49 xor mulr_2_49;
sumr_50<= mulr_1_50 xor mulr_2_50;
sumr_51<= mulr_1_51 xor mulr_2_51;
sumr_52<= mulr_1_52 xor mulr_2_52;
sumr_53<= mulr_1_53 xor mulr_2_53;
sumr_54<= mulr_1_54 xor mulr_2_54;
sumr_55<= mulr_1_55 xor mulr_2_55;
sumr_56<= mulr_1_56 xor mulr_2_56;
sumr_57<= mulr_1_57 xor mulr_2_57;
sumr_58<= mulr_1_58 xor mulr_2_58;
sumr_59<= mulr_1_59 xor mulr_2_59;
sumr_60<= mulr_1_60 xor mulr_2_60;
sumr_61<= mulr_1_61 xor mulr_2_61;
sumr_62<= mulr_1_62 xor mulr_2_62;
sumr_63<= mulr_1_63 xor mulr_2_63;
sumr_64<= mulr_1_64 xor mulr_2_64;
sumr_65<= mulr_1_65 xor mulr_2_65;
sumr_66<= mulr_1_66 xor mulr_2_66;
sumr_67<= mulr_1_67 xor mulr_2_67;
sumr_68<= mulr_1_68 xor mulr_2_68;
sumr_69<= mulr_1_69 xor mulr_2_69;
sumr_70<= mulr_1_70 xor mulr_2_70;
sumr_71<= mulr_1_71 xor mulr_2_71;
sumr_72<= mulr_1_72 xor mulr_2_72;
sumr_73<= mulr_1_73 xor mulr_2_73;
sumr_74<= mulr_1_74 xor mulr_2_74;
sumr_75<= mulr_1_75 xor mulr_2_75;
sumr_76<= mulr_1_76 xor mulr_2_76;
sumr_77<= mulr_1_77 xor mulr_2_77;
sumr_78<= mulr_1_78 xor mulr_2_78;
sumr_79<= mulr_1_79 xor mulr_2_79;
sumr_80<= mulr_1_80 xor mulr_2_80;
sumr_81<= mulr_1_81 xor mulr_2_81;
sumr_82<= mulr_1_82 xor mulr_2_82;
sumr_83<= mulr_1_83 xor mulr_2_83;
sumr_84<= mulr_1_84 xor mulr_2_84;
sumr_85<= mulr_1_85 xor mulr_2_85;
sumr_86<= mulr_1_86 xor mulr_2_86;
sumr_87<= mulr_1_87 xor mulr_2_87;
sumr_88<= mulr_1_88 xor mulr_2_88;
sumr_89<= mulr_1_89 xor mulr_2_89;
sumr_90<= mulr_1_90 xor mulr_2_90;
sumr_91<= mulr_1_91 xor mulr_2_91;
sumr_92<= mulr_1_92 xor mulr_2_92;
sumr_93<= mulr_1_93 xor mulr_2_93;
sumr_94<= mulr_1_94 xor mulr_2_94;
sumr_95<= mulr_1_95 xor mulr_2_95;
sumr_96<= mulr_1_96 xor mulr_2_96;
sumr_97<= mulr_1_97 xor mulr_2_97;
sumr_98<= mulr_1_98 xor mulr_2_98;
sumr_99<= mulr_1_99 xor mulr_2_99;
sumr_100<= mulr_1_100 xor mulr_2_100;
sumr_101<= mulr_1_101 xor mulr_2_101;
sumr_102<= mulr_1_102 xor mulr_2_102;
sumr_103<= mulr_1_103 xor mulr_2_103;
sumr_104<= mulr_1_104 xor mulr_2_104;
sumr_105<= mulr_1_105 xor mulr_2_105;
sumr_106<= mulr_1_106 xor mulr_2_106;
sumr_107<= mulr_1_107 xor mulr_2_107;
sumr_108<= mulr_1_108 xor mulr_2_108;
sumr_109<= mulr_1_109 xor mulr_2_109;
sumr_110<= mulr_1_110 xor mulr_2_110;
sumr_111<= mulr_1_111 xor mulr_2_111;
sumr_112<= mulr_1_112 xor mulr_2_112;
sumr_113<= mulr_1_113 xor mulr_2_113;
sumr_114<= mulr_1_114 xor mulr_2_114;
sumr_115<= mulr_1_115 xor mulr_2_115;
sumr_116<= mulr_1_116 xor mulr_2_116;
sumr_117<= mulr_1_117 xor mulr_2_117;
sumr_118<= mulr_1_118 xor mulr_2_118;
sumr_119<= mulr_1_119 xor mulr_2_119;
sumr_120<= mulr_1_120 xor mulr_2_120;
sumr_121<= mulr_1_121 xor mulr_2_121;
sumr_122<= mulr_1_122 xor mulr_2_122;
sumr_123<= mulr_1_123 xor mulr_2_123;
sumr_124<= mulr_1_124 xor mulr_2_124;
sumr_125<= mulr_1_125 xor mulr_2_125;
sumr_126<= mulr_1_126 xor mulr_2_126;
sumr_127<= mulr_1_127 xor mulr_2_127;
E(126)<=not ( sumr_1(0) or sumr_1(1) or sumr_1(2) or sumr_1(3) or sumr_1(4) or sumr_1(5) or sumr_1(6));
E(125)<=not ( sumr_2(0) or sumr_2(1) or sumr_2(2) or sumr_2(3) or sumr_2(4) or sumr_2(5) or sumr_2(6));
E(124)<=not ( sumr_3(0) or sumr_3(1) or sumr_3(2) or sumr_3(3) or sumr_3(4) or sumr_3(5) or sumr_3(6));
E(123)<=not ( sumr_4(0) or sumr_4(1) or sumr_4(2) or sumr_4(3) or sumr_4(4) or sumr_4(5) or sumr_4(6));
E(122)<=not ( sumr_5(0) or sumr_5(1) or sumr_5(2) or sumr_5(3) or sumr_5(4) or sumr_5(5) or sumr_5(6));
E(121)<=not ( sumr_6(0) or sumr_6(1) or sumr_6(2) or sumr_6(3) or sumr_6(4) or sumr_6(5) or sumr_6(6));
E(120)<=not ( sumr_7(0) or sumr_7(1) or sumr_7(2) or sumr_7(3) or sumr_7(4) or sumr_7(5) or sumr_7(6));
E(119)<=not ( sumr_8(0) or sumr_8(1) or sumr_8(2) or sumr_8(3) or sumr_8(4) or sumr_8(5) or sumr_8(6));
E(118)<=not ( sumr_9(0) or sumr_9(1) or sumr_9(2) or sumr_9(3) or sumr_9(4) or sumr_9(5) or sumr_9(6));
E(117)<=not ( sumr_10(0) or sumr_10(1) or sumr_10(2) or sumr_10(3) or sumr_10(4) or sumr_10(5) or sumr_10(6));
E(116)<=not ( sumr_11(0) or sumr_11(1) or sumr_11(2) or sumr_11(3) or sumr_11(4) or sumr_11(5) or sumr_11(6));
E(115)<=not ( sumr_12(0) or sumr_12(1) or sumr_12(2) or sumr_12(3) or sumr_12(4) or sumr_12(5) or sumr_12(6));
E(114)<=not ( sumr_13(0) or sumr_13(1) or sumr_13(2) or sumr_13(3) or sumr_13(4) or sumr_13(5) or sumr_13(6));
E(113)<=not ( sumr_14(0) or sumr_14(1) or sumr_14(2) or sumr_14(3) or sumr_14(4) or sumr_14(5) or sumr_14(6));
E(112)<=not ( sumr_15(0) or sumr_15(1) or sumr_15(2) or sumr_15(3) or sumr_15(4) or sumr_15(5) or sumr_15(6));
E(111)<=not ( sumr_16(0) or sumr_16(1) or sumr_16(2) or sumr_16(3) or sumr_16(4) or sumr_16(5) or sumr_16(6));
E(110)<=not ( sumr_17(0) or sumr_17(1) or sumr_17(2) or sumr_17(3) or sumr_17(4) or sumr_17(5) or sumr_17(6));
E(109)<=not ( sumr_18(0) or sumr_18(1) or sumr_18(2) or sumr_18(3) or sumr_18(4) or sumr_18(5) or sumr_18(6));
E(108)<=not ( sumr_19(0) or sumr_19(1) or sumr_19(2) or sumr_19(3) or sumr_19(4) or sumr_19(5) or sumr_19(6));
E(107)<=not ( sumr_20(0) or sumr_20(1) or sumr_20(2) or sumr_20(3) or sumr_20(4) or sumr_20(5) or sumr_20(6));
E(106)<=not ( sumr_21(0) or sumr_21(1) or sumr_21(2) or sumr_21(3) or sumr_21(4) or sumr_21(5) or sumr_21(6));
E(105)<=not ( sumr_22(0) or sumr_22(1) or sumr_22(2) or sumr_22(3) or sumr_22(4) or sumr_22(5) or sumr_22(6));
E(104)<=not ( sumr_23(0) or sumr_23(1) or sumr_23(2) or sumr_23(3) or sumr_23(4) or sumr_23(5) or sumr_23(6));
E(103)<=not ( sumr_24(0) or sumr_24(1) or sumr_24(2) or sumr_24(3) or sumr_24(4) or sumr_24(5) or sumr_24(6));
E(102)<=not ( sumr_25(0) or sumr_25(1) or sumr_25(2) or sumr_25(3) or sumr_25(4) or sumr_25(5) or sumr_25(6));
E(101)<=not ( sumr_26(0) or sumr_26(1) or sumr_26(2) or sumr_26(3) or sumr_26(4) or sumr_26(5) or sumr_26(6));
E(100)<=not ( sumr_27(0) or sumr_27(1) or sumr_27(2) or sumr_27(3) or sumr_27(4) or sumr_27(5) or sumr_27(6));
E(99)<=not ( sumr_28(0) or sumr_28(1) or sumr_28(2) or sumr_28(3) or sumr_28(4) or sumr_28(5) or sumr_28(6));
E(98)<=not ( sumr_29(0) or sumr_29(1) or sumr_29(2) or sumr_29(3) or sumr_29(4) or sumr_29(5) or sumr_29(6));
E(97)<=not ( sumr_30(0) or sumr_30(1) or sumr_30(2) or sumr_30(3) or sumr_30(4) or sumr_30(5) or sumr_30(6));
E(96)<=not ( sumr_31(0) or sumr_31(1) or sumr_31(2) or sumr_31(3) or sumr_31(4) or sumr_31(5) or sumr_31(6));
E(95)<=not ( sumr_32(0) or sumr_32(1) or sumr_32(2) or sumr_32(3) or sumr_32(4) or sumr_32(5) or sumr_32(6));
E(94)<=not ( sumr_33(0) or sumr_33(1) or sumr_33(2) or sumr_33(3) or sumr_33(4) or sumr_33(5) or sumr_33(6));
E(93)<=not ( sumr_34(0) or sumr_34(1) or sumr_34(2) or sumr_34(3) or sumr_34(4) or sumr_34(5) or sumr_34(6));
E(92)<=not ( sumr_35(0) or sumr_35(1) or sumr_35(2) or sumr_35(3) or sumr_35(4) or sumr_35(5) or sumr_35(6));
E(91)<=not ( sumr_36(0) or sumr_36(1) or sumr_36(2) or sumr_36(3) or sumr_36(4) or sumr_36(5) or sumr_36(6));
E(90)<=not ( sumr_37(0) or sumr_37(1) or sumr_37(2) or sumr_37(3) or sumr_37(4) or sumr_37(5) or sumr_37(6));
E(89)<=not ( sumr_38(0) or sumr_38(1) or sumr_38(2) or sumr_38(3) or sumr_38(4) or sumr_38(5) or sumr_38(6));
E(88)<=not ( sumr_39(0) or sumr_39(1) or sumr_39(2) or sumr_39(3) or sumr_39(4) or sumr_39(5) or sumr_39(6));
E(87)<=not ( sumr_40(0) or sumr_40(1) or sumr_40(2) or sumr_40(3) or sumr_40(4) or sumr_40(5) or sumr_40(6));
E(86)<=not ( sumr_41(0) or sumr_41(1) or sumr_41(2) or sumr_41(3) or sumr_41(4) or sumr_41(5) or sumr_41(6));
E(85)<=not ( sumr_42(0) or sumr_42(1) or sumr_42(2) or sumr_42(3) or sumr_42(4) or sumr_42(5) or sumr_42(6));
E(84)<=not ( sumr_43(0) or sumr_43(1) or sumr_43(2) or sumr_43(3) or sumr_43(4) or sumr_43(5) or sumr_43(6));
E(83)<=not ( sumr_44(0) or sumr_44(1) or sumr_44(2) or sumr_44(3) or sumr_44(4) or sumr_44(5) or sumr_44(6));
E(82)<=not ( sumr_45(0) or sumr_45(1) or sumr_45(2) or sumr_45(3) or sumr_45(4) or sumr_45(5) or sumr_45(6));
E(81)<=not ( sumr_46(0) or sumr_46(1) or sumr_46(2) or sumr_46(3) or sumr_46(4) or sumr_46(5) or sumr_46(6));
E(80)<=not ( sumr_47(0) or sumr_47(1) or sumr_47(2) or sumr_47(3) or sumr_47(4) or sumr_47(5) or sumr_47(6));
E(79)<=not ( sumr_48(0) or sumr_48(1) or sumr_48(2) or sumr_48(3) or sumr_48(4) or sumr_48(5) or sumr_48(6));
E(78)<=not ( sumr_49(0) or sumr_49(1) or sumr_49(2) or sumr_49(3) or sumr_49(4) or sumr_49(5) or sumr_49(6));
E(77)<=not ( sumr_50(0) or sumr_50(1) or sumr_50(2) or sumr_50(3) or sumr_50(4) or sumr_50(5) or sumr_50(6));
E(76)<=not ( sumr_51(0) or sumr_51(1) or sumr_51(2) or sumr_51(3) or sumr_51(4) or sumr_51(5) or sumr_51(6));
E(75)<=not ( sumr_52(0) or sumr_52(1) or sumr_52(2) or sumr_52(3) or sumr_52(4) or sumr_52(5) or sumr_52(6));
E(74)<=not ( sumr_53(0) or sumr_53(1) or sumr_53(2) or sumr_53(3) or sumr_53(4) or sumr_53(5) or sumr_53(6));
E(73)<=not ( sumr_54(0) or sumr_54(1) or sumr_54(2) or sumr_54(3) or sumr_54(4) or sumr_54(5) or sumr_54(6));
E(72)<=not ( sumr_55(0) or sumr_55(1) or sumr_55(2) or sumr_55(3) or sumr_55(4) or sumr_55(5) or sumr_55(6));
E(71)<=not ( sumr_56(0) or sumr_56(1) or sumr_56(2) or sumr_56(3) or sumr_56(4) or sumr_56(5) or sumr_56(6));
E(70)<=not ( sumr_57(0) or sumr_57(1) or sumr_57(2) or sumr_57(3) or sumr_57(4) or sumr_57(5) or sumr_57(6));
E(69)<=not ( sumr_58(0) or sumr_58(1) or sumr_58(2) or sumr_58(3) or sumr_58(4) or sumr_58(5) or sumr_58(6));
E(68)<=not ( sumr_59(0) or sumr_59(1) or sumr_59(2) or sumr_59(3) or sumr_59(4) or sumr_59(5) or sumr_59(6));
E(67)<=not ( sumr_60(0) or sumr_60(1) or sumr_60(2) or sumr_60(3) or sumr_60(4) or sumr_60(5) or sumr_60(6));
E(66)<=not ( sumr_61(0) or sumr_61(1) or sumr_61(2) or sumr_61(3) or sumr_61(4) or sumr_61(5) or sumr_61(6));
E(65)<=not ( sumr_62(0) or sumr_62(1) or sumr_62(2) or sumr_62(3) or sumr_62(4) or sumr_62(5) or sumr_62(6));
E(64)<=not ( sumr_63(0) or sumr_63(1) or sumr_63(2) or sumr_63(3) or sumr_63(4) or sumr_63(5) or sumr_63(6));
E(63)<=not ( sumr_64(0) or sumr_64(1) or sumr_64(2) or sumr_64(3) or sumr_64(4) or sumr_64(5) or sumr_64(6));
E(62)<=not ( sumr_65(0) or sumr_65(1) or sumr_65(2) or sumr_65(3) or sumr_65(4) or sumr_65(5) or sumr_65(6));
E(61)<=not ( sumr_66(0) or sumr_66(1) or sumr_66(2) or sumr_66(3) or sumr_66(4) or sumr_66(5) or sumr_66(6));
E(60)<=not ( sumr_67(0) or sumr_67(1) or sumr_67(2) or sumr_67(3) or sumr_67(4) or sumr_67(5) or sumr_67(6));
E(59)<=not ( sumr_68(0) or sumr_68(1) or sumr_68(2) or sumr_68(3) or sumr_68(4) or sumr_68(5) or sumr_68(6));
E(58)<=not ( sumr_69(0) or sumr_69(1) or sumr_69(2) or sumr_69(3) or sumr_69(4) or sumr_69(5) or sumr_69(6));
E(57)<=not ( sumr_70(0) or sumr_70(1) or sumr_70(2) or sumr_70(3) or sumr_70(4) or sumr_70(5) or sumr_70(6));
E(56)<=not ( sumr_71(0) or sumr_71(1) or sumr_71(2) or sumr_71(3) or sumr_71(4) or sumr_71(5) or sumr_71(6));
E(55)<=not ( sumr_72(0) or sumr_72(1) or sumr_72(2) or sumr_72(3) or sumr_72(4) or sumr_72(5) or sumr_72(6));
E(54)<=not ( sumr_73(0) or sumr_73(1) or sumr_73(2) or sumr_73(3) or sumr_73(4) or sumr_73(5) or sumr_73(6));
E(53)<=not ( sumr_74(0) or sumr_74(1) or sumr_74(2) or sumr_74(3) or sumr_74(4) or sumr_74(5) or sumr_74(6));
E(52)<=not ( sumr_75(0) or sumr_75(1) or sumr_75(2) or sumr_75(3) or sumr_75(4) or sumr_75(5) or sumr_75(6));
E(51)<=not ( sumr_76(0) or sumr_76(1) or sumr_76(2) or sumr_76(3) or sumr_76(4) or sumr_76(5) or sumr_76(6));
E(50)<=not ( sumr_77(0) or sumr_77(1) or sumr_77(2) or sumr_77(3) or sumr_77(4) or sumr_77(5) or sumr_77(6));
E(49)<=not ( sumr_78(0) or sumr_78(1) or sumr_78(2) or sumr_78(3) or sumr_78(4) or sumr_78(5) or sumr_78(6));
E(48)<=not ( sumr_79(0) or sumr_79(1) or sumr_79(2) or sumr_79(3) or sumr_79(4) or sumr_79(5) or sumr_79(6));
E(47)<=not ( sumr_80(0) or sumr_80(1) or sumr_80(2) or sumr_80(3) or sumr_80(4) or sumr_80(5) or sumr_80(6));
E(46)<=not ( sumr_81(0) or sumr_81(1) or sumr_81(2) or sumr_81(3) or sumr_81(4) or sumr_81(5) or sumr_81(6));
E(45)<=not ( sumr_82(0) or sumr_82(1) or sumr_82(2) or sumr_82(3) or sumr_82(4) or sumr_82(5) or sumr_82(6));
E(44)<=not ( sumr_83(0) or sumr_83(1) or sumr_83(2) or sumr_83(3) or sumr_83(4) or sumr_83(5) or sumr_83(6));
E(43)<=not ( sumr_84(0) or sumr_84(1) or sumr_84(2) or sumr_84(3) or sumr_84(4) or sumr_84(5) or sumr_84(6));
E(42)<=not ( sumr_85(0) or sumr_85(1) or sumr_85(2) or sumr_85(3) or sumr_85(4) or sumr_85(5) or sumr_85(6));
E(41)<=not ( sumr_86(0) or sumr_86(1) or sumr_86(2) or sumr_86(3) or sumr_86(4) or sumr_86(5) or sumr_86(6));
E(40)<=not ( sumr_87(0) or sumr_87(1) or sumr_87(2) or sumr_87(3) or sumr_87(4) or sumr_87(5) or sumr_87(6));
E(39)<=not ( sumr_88(0) or sumr_88(1) or sumr_88(2) or sumr_88(3) or sumr_88(4) or sumr_88(5) or sumr_88(6));
E(38)<=not ( sumr_89(0) or sumr_89(1) or sumr_89(2) or sumr_89(3) or sumr_89(4) or sumr_89(5) or sumr_89(6));
E(37)<=not ( sumr_90(0) or sumr_90(1) or sumr_90(2) or sumr_90(3) or sumr_90(4) or sumr_90(5) or sumr_90(6));
E(36)<=not ( sumr_91(0) or sumr_91(1) or sumr_91(2) or sumr_91(3) or sumr_91(4) or sumr_91(5) or sumr_91(6));
E(35)<=not ( sumr_92(0) or sumr_92(1) or sumr_92(2) or sumr_92(3) or sumr_92(4) or sumr_92(5) or sumr_92(6));
E(34)<=not ( sumr_93(0) or sumr_93(1) or sumr_93(2) or sumr_93(3) or sumr_93(4) or sumr_93(5) or sumr_93(6));
E(33)<=not ( sumr_94(0) or sumr_94(1) or sumr_94(2) or sumr_94(3) or sumr_94(4) or sumr_94(5) or sumr_94(6));
E(32)<=not ( sumr_95(0) or sumr_95(1) or sumr_95(2) or sumr_95(3) or sumr_95(4) or sumr_95(5) or sumr_95(6));
E(31)<=not ( sumr_96(0) or sumr_96(1) or sumr_96(2) or sumr_96(3) or sumr_96(4) or sumr_96(5) or sumr_96(6));
E(30)<=not ( sumr_97(0) or sumr_97(1) or sumr_97(2) or sumr_97(3) or sumr_97(4) or sumr_97(5) or sumr_97(6));
E(29)<=not ( sumr_98(0) or sumr_98(1) or sumr_98(2) or sumr_98(3) or sumr_98(4) or sumr_98(5) or sumr_98(6));
E(28)<=not ( sumr_99(0) or sumr_99(1) or sumr_99(2) or sumr_99(3) or sumr_99(4) or sumr_99(5) or sumr_99(6));
E(27)<=not ( sumr_100(0) or sumr_100(1) or sumr_100(2) or sumr_100(3) or sumr_100(4) or sumr_100(5) or sumr_100(6));
E(26)<=not ( sumr_101(0) or sumr_101(1) or sumr_101(2) or sumr_101(3) or sumr_101(4) or sumr_101(5) or sumr_101(6));
E(25)<=not ( sumr_102(0) or sumr_102(1) or sumr_102(2) or sumr_102(3) or sumr_102(4) or sumr_102(5) or sumr_102(6));
E(24)<=not ( sumr_103(0) or sumr_103(1) or sumr_103(2) or sumr_103(3) or sumr_103(4) or sumr_103(5) or sumr_103(6));
E(23)<=not ( sumr_104(0) or sumr_104(1) or sumr_104(2) or sumr_104(3) or sumr_104(4) or sumr_104(5) or sumr_104(6));
E(22)<=not ( sumr_105(0) or sumr_105(1) or sumr_105(2) or sumr_105(3) or sumr_105(4) or sumr_105(5) or sumr_105(6));
E(21)<=not ( sumr_106(0) or sumr_106(1) or sumr_106(2) or sumr_106(3) or sumr_106(4) or sumr_106(5) or sumr_106(6));
E(20)<=not ( sumr_107(0) or sumr_107(1) or sumr_107(2) or sumr_107(3) or sumr_107(4) or sumr_107(5) or sumr_107(6));
E(19)<=not ( sumr_108(0) or sumr_108(1) or sumr_108(2) or sumr_108(3) or sumr_108(4) or sumr_108(5) or sumr_108(6));
E(18)<=not ( sumr_109(0) or sumr_109(1) or sumr_109(2) or sumr_109(3) or sumr_109(4) or sumr_109(5) or sumr_109(6));
E(17)<=not ( sumr_110(0) or sumr_110(1) or sumr_110(2) or sumr_110(3) or sumr_110(4) or sumr_110(5) or sumr_110(6));
E(16)<=not ( sumr_111(0) or sumr_111(1) or sumr_111(2) or sumr_111(3) or sumr_111(4) or sumr_111(5) or sumr_111(6));
E(15)<=not ( sumr_112(0) or sumr_112(1) or sumr_112(2) or sumr_112(3) or sumr_112(4) or sumr_112(5) or sumr_112(6));
E(14)<=not ( sumr_113(0) or sumr_113(1) or sumr_113(2) or sumr_113(3) or sumr_113(4) or sumr_113(5) or sumr_113(6));
E(13)<=not ( sumr_114(0) or sumr_114(1) or sumr_114(2) or sumr_114(3) or sumr_114(4) or sumr_114(5) or sumr_114(6));
E(12)<=not ( sumr_115(0) or sumr_115(1) or sumr_115(2) or sumr_115(3) or sumr_115(4) or sumr_115(5) or sumr_115(6));
E(11)<=not ( sumr_116(0) or sumr_116(1) or sumr_116(2) or sumr_116(3) or sumr_116(4) or sumr_116(5) or sumr_116(6));
E(10)<=not ( sumr_117(0) or sumr_117(1) or sumr_117(2) or sumr_117(3) or sumr_117(4) or sumr_117(5) or sumr_117(6));
E(9)<=not ( sumr_118(0) or sumr_118(1) or sumr_118(2) or sumr_118(3) or sumr_118(4) or sumr_118(5) or sumr_118(6));
E(8)<=not ( sumr_119(0) or sumr_119(1) or sumr_119(2) or sumr_119(3) or sumr_119(4) or sumr_119(5) or sumr_119(6));
E(7)<=not ( sumr_120(0) or sumr_120(1) or sumr_120(2) or sumr_120(3) or sumr_120(4) or sumr_120(5) or sumr_120(6));
E(6)<=not ( sumr_121(0) or sumr_121(1) or sumr_121(2) or sumr_121(3) or sumr_121(4) or sumr_121(5) or sumr_121(6));
E(5)<=not ( sumr_122(0) or sumr_122(1) or sumr_122(2) or sumr_122(3) or sumr_122(4) or sumr_122(5) or sumr_122(6));
E(4)<=not ( sumr_123(0) or sumr_123(1) or sumr_123(2) or sumr_123(3) or sumr_123(4) or sumr_123(5) or sumr_123(6));
E(3)<=not ( sumr_124(0) or sumr_124(1) or sumr_124(2) or sumr_124(3) or sumr_124(4) or sumr_124(5) or sumr_124(6));
E(2)<=not ( sumr_125(0) or sumr_125(1) or sumr_125(2) or sumr_125(3) or sumr_125(4) or sumr_125(5) or sumr_125(6));
E(1)<=not ( sumr_126(0) or sumr_126(1) or sumr_126(2) or sumr_126(3) or sumr_126(4) or sumr_126(5) or sumr_126(6));
E(0)<=not ( sumr_127(0) or sumr_127(1) or sumr_127(2) or sumr_127(3) or sumr_127(4) or sumr_127(5) or sumr_127(6));
end arch;
