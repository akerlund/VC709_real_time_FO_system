library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.ALL;
package word_expander_package_for_D64_N99 is

    constant INPUT_WIDTH : integer := 64;
    constant OUTPUT_WIDTH : integer := 99;
    constant INPUT_ROM_ROWS : integer := 16;


    type ROM_type_expanded is array (0 to (INPUT_WIDTH*INPUT_ROM_ROWS-1)) of std_logic_vector((OUTPUT_WIDTH-1) downto 0);
    constant ROM_expanded : ROM_type_expanded := (
            "000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000",
            "111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
            "000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000",
            "111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111",
            "000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000",
            "011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000",
            "111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
            "000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000",
            "111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111",
            "000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
            "111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111",
            "000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000",
            "111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
            "000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000",
            "111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111",
            "000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000",
            "000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000",
            "111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111",
            "000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000",
            "111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111",
            "000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000",
            "111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111",
            "000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000",
            "111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111",
            "000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000",
            "111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111",
            "000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110",
            "000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000",
            "111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111",
            "000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000",
            "111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111",
            "000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000",
            "111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111",
            "000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000",
            "111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111",
            "000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000",
            "111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111",
            "100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111",
            "000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000",
            "111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111",
            "000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
            "111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111",
            "000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000",
            "111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111",
            "000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000",
            "111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111",
            "000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000",
            "111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111",
            "111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111",
            "000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000",
            "111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111",
            "000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
            "111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111",
            "000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000",
            "111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111",
            "000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000",
            "111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111",
            "000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000",
            "111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001",
            "111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
            "000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000",
            "111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111",
            "000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
            "111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111",
            "000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000",
            "111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
            "000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000",
            "111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111",
            "000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000",
            "011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000",
            "111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
            "000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000",
            "111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111",
            "000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
            "111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111",
            "000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000",
            "111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
            "000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000",
            "111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111",
            "000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000",
            "000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000",
            "111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111",
            "000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000",
            "111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111",
            "000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000",
            "111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111",
            "000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000",
            "111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111",
            "000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000",
            "111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111",
            "000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110",
            "000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000",
            "111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111",
            "000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000",
            "111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111",
            "000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000",
            "111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111",
            "000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000",
            "111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111",
            "000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000",
            "111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111",
            "100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111",
            "000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000",
            "111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111",
            "000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
            "111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111",
            "000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000",
            "111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111",
            "000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000",
            "111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111",
            "000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000",
            "111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111",
            "111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111",
            "000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000",
            "111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111",
            "000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
            "111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111",
            "000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000",
            "111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111",
            "000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000",
            "111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111",
            "000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000",
            "111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001",
            "111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
            "000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000",
            "111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111",
            "000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
            "111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111",
            "000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000",
            "111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
            "000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000",
            "111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111",
            "000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000",
            "011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000",
            "111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
            "000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000",
            "111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111",
            "000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
            "111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111",
            "000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000",
            "111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
            "000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000",
            "111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111",
            "000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000",
            "000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000",
            "111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111",
            "000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000",
            "111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111",
            "000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000",
            "111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111",
            "000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000",
            "111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111",
            "000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000",
            "111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111",
            "000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110",
            "000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000",
            "111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111",
            "000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000",
            "111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111",
            "000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000",
            "111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111",
            "000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000",
            "111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111",
            "000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000",
            "111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111",
            "100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111",
            "000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000",
            "111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111",
            "000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
            "111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111",
            "000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000",
            "111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111",
            "000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000",
            "111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111",
            "000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000",
            "111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111",
            "111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111",
            "000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000",
            "111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111",
            "000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
            "111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111",
            "000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000",
            "111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111",
            "000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000",
            "111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111",
            "000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000",
            "111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001",
            "111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
            "000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000",
            "111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111",
            "000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
            "111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111",
            "000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000",
            "111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
            "000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000",
            "111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111",
            "000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000",
            "011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000",
            "111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
            "000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000",
            "111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111",
            "000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
            "111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111",
            "000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000",
            "111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
            "000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000",
            "111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111",
            "000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000",
            "000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000",
            "111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111",
            "000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000",
            "111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111",
            "000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000",
            "111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111",
            "000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000",
            "111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111",
            "000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000",
            "111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111",
            "000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110",
            "000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000",
            "111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111",
            "000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000",
            "111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111",
            "000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000",
            "111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111",
            "000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000",
            "111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111",
            "000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000",
            "111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111",
            "100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111",
            "000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000",
            "111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111",
            "000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
            "111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111",
            "000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000",
            "111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111",
            "000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000",
            "111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111",
            "000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000",
            "111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111",
            "111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111",
            "000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000",
            "111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111",
            "000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
            "111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111",
            "000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000",
            "111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111",
            "000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000",
            "111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111",
            "000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000",
            "111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001",
            "111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
            "000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000",
            "111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111",
            "000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
            "111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111",
            "000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000",
            "111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
            "000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000",
            "111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111",
            "000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000",
            "011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000",
            "111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
            "000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000",
            "111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111",
            "000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
            "111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111",
            "000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000",
            "111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
            "000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000",
            "111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111",
            "000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000",
            "000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000",
            "111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111",
            "000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000",
            "111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111",
            "000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000",
            "111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111",
            "000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000",
            "111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111",
            "000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000",
            "111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111",
            "000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110",
            "000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000",
            "111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111",
            "000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000",
            "111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111",
            "000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000",
            "111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111",
            "000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000",
            "111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111",
            "000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000",
            "111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111",
            "100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111",
            "000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000",
            "111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111",
            "000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
            "111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111",
            "000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000",
            "111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111",
            "000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000",
            "111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111",
            "000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000",
            "111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111",
            "111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111",
            "000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000",
            "111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111",
            "000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
            "111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111",
            "000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000",
            "111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111",
            "000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000",
            "111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111",
            "000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000",
            "111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001",
            "111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
            "000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000",
            "111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111",
            "000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
            "111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111",
            "000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000",
            "111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
            "000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000",
            "111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111",
            "000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000",
            "011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000",
            "111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
            "000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000",
            "111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111",
            "000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
            "111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111",
            "000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000",
            "111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
            "000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000",
            "111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111",
            "000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000",
            "000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000",
            "111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111",
            "000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000",
            "111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111",
            "000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000",
            "111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111",
            "000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000",
            "111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111",
            "000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000",
            "111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111",
            "000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110",
            "000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000",
            "111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111",
            "000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000",
            "111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111",
            "000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000",
            "111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111",
            "000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000",
            "111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111",
            "000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000",
            "111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111",
            "100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111",
            "000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000",
            "111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111",
            "000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
            "111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111",
            "000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000",
            "111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111",
            "000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000",
            "111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111",
            "000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000",
            "111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111",
            "111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111",
            "000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000",
            "111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111",
            "000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
            "111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111",
            "000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000",
            "111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111",
            "000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000",
            "111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111",
            "000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000",
            "111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001",
            "111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
            "000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000",
            "111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111",
            "000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
            "111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111",
            "000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000",
            "111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
            "000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000",
            "111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111",
            "000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000",
            "011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000",
            "111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
            "000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000",
            "111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111",
            "000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
            "111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111",
            "000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000",
            "111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
            "000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000",
            "111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111",
            "000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000",
            "000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000",
            "111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111",
            "000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000",
            "111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111",
            "000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000",
            "111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111",
            "000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000",
            "111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111",
            "000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000",
            "111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111",
            "000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110",
            "000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000",
            "111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111",
            "000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000",
            "111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111",
            "000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000",
            "111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111",
            "000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000",
            "111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111",
            "000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000",
            "111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111",
            "100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111",
            "000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000",
            "111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111",
            "000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
            "111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111",
            "000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000",
            "111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111",
            "000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000",
            "111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111",
            "000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000",
            "111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111",
            "111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111",
            "000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000",
            "111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111",
            "000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
            "111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111",
            "000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000",
            "111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111",
            "000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000",
            "111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111",
            "000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000",
            "111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001",
            "111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
            "000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000",
            "111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111",
            "000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
            "111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111",
            "000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000",
            "111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
            "000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000",
            "111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111",
            "000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000",
            "011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000",
            "111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
            "000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000",
            "111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111",
            "000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
            "111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111",
            "000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000",
            "111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
            "000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000",
            "111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111",
            "000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000",
            "000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000",
            "111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111",
            "000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000",
            "111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111",
            "000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000",
            "111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111",
            "000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000",
            "111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111",
            "000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000",
            "111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111",
            "000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110",
            "000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000",
            "111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111",
            "000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000",
            "111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111",
            "000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000",
            "111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111",
            "000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000",
            "111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111",
            "000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000",
            "111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111",
            "100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111",
            "000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000",
            "111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111",
            "000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
            "111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111",
            "000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000",
            "111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111",
            "000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000",
            "111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111",
            "000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000",
            "111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111",
            "111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111",
            "000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000",
            "111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111",
            "000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
            "111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111",
            "000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000",
            "111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111",
            "000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000",
            "111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111",
            "000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000",
            "111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001",
            "111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
            "000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000",
            "111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111",
            "000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
            "111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111"
    );

    type ROM_type_data is array (0 to (INPUT_ROM_ROWS-1)) of std_logic_vector((INPUT_WIDTH-1) downto 0);
    constant ROM_data : ROM_type_data := (
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000"
    );

    function ROM_send_data(index : integer) return std_logic_vector;    function ROM_D64_N99(index : integer) return std_logic_vector;

end word_expander_package_for_D64_N99;

package body word_expander_package_for_D64_N99 is

    function ROM_send_data(index : integer) return std_logic_vector is
    begin
        return ROM_data(index);
    end ROM_send_data;


    function ROM_D64_N99(index : integer) return std_logic_vector is
    begin
        return ROM_expanded(index);
    end ROM_D64_N99;


end word_expander_package_for_D64_N99;