library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.ALL;
package word_expander_package_for_D64_N106 is

    constant INPUT_WIDTH : integer := 64;
    constant OUTPUT_WIDTH : integer := 106;
    constant INPUT_ROM_ROWS : integer := 16;


    type ROM_type_expanded is array (0 to (INPUT_WIDTH*INPUT_ROM_ROWS-1)) of std_logic_vector((OUTPUT_WIDTH-1) downto 0);
    constant ROM_expanded : ROM_type_expanded := (
            "0000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "1111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "0000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "1111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "0000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "1111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "0000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "1111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "0000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "1100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "0000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "0000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "1111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "0000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "1111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "0000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "1111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "0011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "1111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "0000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "1111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "0000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "1111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "0000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "1111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "0000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "1100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "0000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "0000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "1111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "0000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "1111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "0000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "1111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "0011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "1111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "0000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "1111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "0000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "1111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "0000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "1111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "0000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "1100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "0000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "0000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "1111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "0000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "1111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "0000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "1111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "0011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "1111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "0000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "1111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "0000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "1111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "0000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "1111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "0000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "1100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "0000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "0000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "1111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "0000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "1111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "0000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "1111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "0011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "1111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "0000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "1111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "0000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "1111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "0000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "1111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "0000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "1100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "0000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "0000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "1111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "0000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "1111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "0000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "1111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "0011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "1111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "0000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "1111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "0000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "1111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "0000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "1111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "0000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "1100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "0000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "0000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "1111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "0000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "1111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "0000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "1111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "0011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "1111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "0000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "1111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "0000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "1111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "0000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "1111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "0000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "1100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "0000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "0000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "1111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "0000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "1111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "0000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "1111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "0011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "1111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "0000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "1111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "0000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "1111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "0000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "1111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "0000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "1100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "0000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "0000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "1111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "0000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "1111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "0000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "1111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "0011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "1111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "0000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "1111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "0000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "1111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "0000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "1111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "0000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "1100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "0000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "0000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "1111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "0000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "1111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "0000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "1111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "0011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "1111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "0000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "1111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "0000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "1111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "0000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "1111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "0000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "1100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "0000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "0000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "1111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "0000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "1111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "0000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "1111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "0011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "1111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "0000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "1111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "0000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "1111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "0000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "1111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "0000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "1100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "0000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "0000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "1111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "0000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "1111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "0000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "1111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "0011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "1111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "0000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "1111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "0000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "1111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "0000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "1111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "0000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "1100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "0000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "0000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "1111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "0000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "1111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "0000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "1111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "0011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "1111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "0000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "1111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "0000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "1111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "0000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "1111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "0000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "1100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "0000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "0000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "1111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "0000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "1111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "0000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "1111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "0011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "1111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "0000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "1111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "0000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "1111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "0000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "1111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "0000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "1100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "0000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "0000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "1111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "0000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "1111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "0000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "1111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "0011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "1111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "0000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "1111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "0000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "1111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "0000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "1111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "0000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "1100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "0000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "0000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "1111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "0000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "1111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "0000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "1111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "0011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "1111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "0000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "1111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "0000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "1111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "0000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "1111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "0000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "1100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "0000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "0000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "1111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "0000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "1111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "0000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "1111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "0011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111"
    );

    type ROM_type_data is array (0 to (INPUT_ROM_ROWS-1)) of std_logic_vector((INPUT_WIDTH-1) downto 0);
    constant ROM_data : ROM_type_data := (
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000"
    );

    function ROM_send_data(index : integer) return std_logic_vector;    function ROM_D64_N106(index : integer) return std_logic_vector;

end word_expander_package_for_D64_N106;

package body word_expander_package_for_D64_N106 is

    function ROM_send_data(index : integer) return std_logic_vector is
    begin
        return ROM_data(index);
    end ROM_send_data;


    function ROM_D64_N106(index : integer) return std_logic_vector is
    begin
        return ROM_expanded(index);
    end ROM_D64_N106;


end word_expander_package_for_D64_N106;