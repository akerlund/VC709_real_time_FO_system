----------------------------------------------------------------------------------
    -- Company:  Chalmers
    -- Engineer: Fredrik Åkerlund
    -- 
    -- Create Date: Mon Jul 24 13:30:05 2017

    -- Design Name: 
    -- Module Name: word_expander_64IN_to_1003OUT - arch_word_expander_64IN_to_1003OUT
    -- Project Name: 
    -- Target Devices: 
    -- Tool Versions: 
    -- Description: 
    -- 
    -- Dependencies: 
    -- 
    -- Revision:
    -- Revision 0.01 - File Created
    -- Additional Comments:
    -- 
    ----------------------------------------------------------------------------------


    library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;

    -- Uncomment the following library declaration if using
    -- arithmetic functions with Signed or Unsigned values
    use IEEE.NUMERIC_STD.ALL;

    -- Uncomment the following library declaration if instantiating
    -- any Xilinx leaf cells in this code.
    --library UNISIM;
    --use UNISIM.VComponents.all;
    entity word_expander_64IN_to_1003OUT is

    generic(
        IN_WIDTH  : integer := 64;
        OUT_WIDTH : integer := 1003
    );
    port(
        user_clk  : in  std_logic;       
        reset_in  : in  std_logic;
        enable_in : in  std_logic;

        in_rdy    : in  std_logic;
        data_in   : in  std_logic_vector(IN_WIDTH-1 downto 0);

        buf_out   : out std_logic_vector(OUT_WIDTH-1 downto 0);
        out_rdy   : out std_logic

        );
    end word_expander_64IN_to_1003OUT;
architecture arch_word_expander_64IN_to_1003OUT of word_expander_64IN_to_1003OUT is

        constant BUF_WIDTH : integer := (OUT_WIDTH + IN_WIDTH);

        signal buf_input_r  : std_logic_vector(BUF_WIDTH-1 downto 0);
        signal buf_output_r : std_logic_vector(OUT_WIDTH-1 downto 0);
        signal out_rdy_r    : std_logic;

        signal bits_in_buffer : integer range 0 to BUF_WIDTH;

    begin

    output_reg_process:
    process(reset_in, user_clk, enable_in)
    begin
        if reset_in = '0' then
            buf_out <= (others=>'0');
            out_rdy <= '0';
        elsif rising_edge(user_clk) then
            if enable_in = '1' then
                buf_out <= buf_output_r;
                out_rdy <= out_rdy_r;
            end if;
        end if;
    end process;


    the_buffing_process:
    process(reset_in, user_clk, in_rdy, enable_in)
    begin
        if reset_in = '0' then

            buf_input_r  <= (others=>'0');
            buf_output_r <= (others=>'0');

            bits_in_buffer <= 0;

            out_rdy_r <= '0';

        elsif rising_edge(user_clk) then
            if in_rdy = '1' and enable_in = '1' then
            if bits_in_buffer >= 939 then
                out_rdy_r <= '1';
                case bits_in_buffer is
                    when 939 =>
                        buf_output_r(938 downto 0)   <= buf_input_r(938 downto 0);
                        buf_output_r(1002 downto 939) <= data_in(63 downto 0);
                        buf_input_r                  <= (others=>'0');
                        bits_in_buffer               <= 0;
                    when 940 =>
                        buf_output_r(939 downto 0)   <= buf_input_r(939 downto 0);
                        buf_output_r(1002 downto 940) <= data_in(62 downto 0);
                        buf_input_r (0 downto 0)     <= data_in(63 downto 63);
                        bits_in_buffer               <= 1;
                    when 941 =>
                        buf_output_r(940 downto 0)   <= buf_input_r(940 downto 0);
                        buf_output_r(1002 downto 941) <= data_in(61 downto 0);
                        buf_input_r (1 downto 0)     <= data_in(63 downto 62);
                        bits_in_buffer               <= 2;
                    when 942 =>
                        buf_output_r(941 downto 0)   <= buf_input_r(941 downto 0);
                        buf_output_r(1002 downto 942) <= data_in(60 downto 0);
                        buf_input_r (2 downto 0)     <= data_in(63 downto 61);
                        bits_in_buffer               <= 3;
                    when 943 =>
                        buf_output_r(942 downto 0)   <= buf_input_r(942 downto 0);
                        buf_output_r(1002 downto 943) <= data_in(59 downto 0);
                        buf_input_r (3 downto 0)     <= data_in(63 downto 60);
                        bits_in_buffer               <= 4;
                    when 944 =>
                        buf_output_r(943 downto 0)   <= buf_input_r(943 downto 0);
                        buf_output_r(1002 downto 944) <= data_in(58 downto 0);
                        buf_input_r (4 downto 0)     <= data_in(63 downto 59);
                        bits_in_buffer               <= 5;
                    when 945 =>
                        buf_output_r(944 downto 0)   <= buf_input_r(944 downto 0);
                        buf_output_r(1002 downto 945) <= data_in(57 downto 0);
                        buf_input_r (5 downto 0)     <= data_in(63 downto 58);
                        bits_in_buffer               <= 6;
                    when 946 =>
                        buf_output_r(945 downto 0)   <= buf_input_r(945 downto 0);
                        buf_output_r(1002 downto 946) <= data_in(56 downto 0);
                        buf_input_r (6 downto 0)     <= data_in(63 downto 57);
                        bits_in_buffer               <= 7;
                    when 947 =>
                        buf_output_r(946 downto 0)   <= buf_input_r(946 downto 0);
                        buf_output_r(1002 downto 947) <= data_in(55 downto 0);
                        buf_input_r (7 downto 0)     <= data_in(63 downto 56);
                        bits_in_buffer               <= 8;
                    when 948 =>
                        buf_output_r(947 downto 0)   <= buf_input_r(947 downto 0);
                        buf_output_r(1002 downto 948) <= data_in(54 downto 0);
                        buf_input_r (8 downto 0)     <= data_in(63 downto 55);
                        bits_in_buffer               <= 9;
                    when 949 =>
                        buf_output_r(948 downto 0)   <= buf_input_r(948 downto 0);
                        buf_output_r(1002 downto 949) <= data_in(53 downto 0);
                        buf_input_r (9 downto 0)     <= data_in(63 downto 54);
                        bits_in_buffer               <= 10;
                    when 950 =>
                        buf_output_r(949 downto 0)   <= buf_input_r(949 downto 0);
                        buf_output_r(1002 downto 950) <= data_in(52 downto 0);
                        buf_input_r (10 downto 0)    <= data_in(63 downto 53);
                        bits_in_buffer               <= 11;
                    when 951 =>
                        buf_output_r(950 downto 0)   <= buf_input_r(950 downto 0);
                        buf_output_r(1002 downto 951) <= data_in(51 downto 0);
                        buf_input_r (11 downto 0)    <= data_in(63 downto 52);
                        bits_in_buffer               <= 12;
                    when 952 =>
                        buf_output_r(951 downto 0)   <= buf_input_r(951 downto 0);
                        buf_output_r(1002 downto 952) <= data_in(50 downto 0);
                        buf_input_r (12 downto 0)    <= data_in(63 downto 51);
                        bits_in_buffer               <= 13;
                    when 953 =>
                        buf_output_r(952 downto 0)   <= buf_input_r(952 downto 0);
                        buf_output_r(1002 downto 953) <= data_in(49 downto 0);
                        buf_input_r (13 downto 0)    <= data_in(63 downto 50);
                        bits_in_buffer               <= 14;
                    when 954 =>
                        buf_output_r(953 downto 0)   <= buf_input_r(953 downto 0);
                        buf_output_r(1002 downto 954) <= data_in(48 downto 0);
                        buf_input_r (14 downto 0)    <= data_in(63 downto 49);
                        bits_in_buffer               <= 15;
                    when 955 =>
                        buf_output_r(954 downto 0)   <= buf_input_r(954 downto 0);
                        buf_output_r(1002 downto 955) <= data_in(47 downto 0);
                        buf_input_r (15 downto 0)    <= data_in(63 downto 48);
                        bits_in_buffer               <= 16;
                    when 956 =>
                        buf_output_r(955 downto 0)   <= buf_input_r(955 downto 0);
                        buf_output_r(1002 downto 956) <= data_in(46 downto 0);
                        buf_input_r (16 downto 0)    <= data_in(63 downto 47);
                        bits_in_buffer               <= 17;
                    when 957 =>
                        buf_output_r(956 downto 0)   <= buf_input_r(956 downto 0);
                        buf_output_r(1002 downto 957) <= data_in(45 downto 0);
                        buf_input_r (17 downto 0)    <= data_in(63 downto 46);
                        bits_in_buffer               <= 18;
                    when 958 =>
                        buf_output_r(957 downto 0)   <= buf_input_r(957 downto 0);
                        buf_output_r(1002 downto 958) <= data_in(44 downto 0);
                        buf_input_r (18 downto 0)    <= data_in(63 downto 45);
                        bits_in_buffer               <= 19;
                    when 959 =>
                        buf_output_r(958 downto 0)   <= buf_input_r(958 downto 0);
                        buf_output_r(1002 downto 959) <= data_in(43 downto 0);
                        buf_input_r (19 downto 0)    <= data_in(63 downto 44);
                        bits_in_buffer               <= 20;
                    when 960 =>
                        buf_output_r(959 downto 0)   <= buf_input_r(959 downto 0);
                        buf_output_r(1002 downto 960) <= data_in(42 downto 0);
                        buf_input_r (20 downto 0)    <= data_in(63 downto 43);
                        bits_in_buffer               <= 21;
                    when 961 =>
                        buf_output_r(960 downto 0)   <= buf_input_r(960 downto 0);
                        buf_output_r(1002 downto 961) <= data_in(41 downto 0);
                        buf_input_r (21 downto 0)    <= data_in(63 downto 42);
                        bits_in_buffer               <= 22;
                    when 962 =>
                        buf_output_r(961 downto 0)   <= buf_input_r(961 downto 0);
                        buf_output_r(1002 downto 962) <= data_in(40 downto 0);
                        buf_input_r (22 downto 0)    <= data_in(63 downto 41);
                        bits_in_buffer               <= 23;
                    when 963 =>
                        buf_output_r(962 downto 0)   <= buf_input_r(962 downto 0);
                        buf_output_r(1002 downto 963) <= data_in(39 downto 0);
                        buf_input_r (23 downto 0)    <= data_in(63 downto 40);
                        bits_in_buffer               <= 24;
                    when 964 =>
                        buf_output_r(963 downto 0)   <= buf_input_r(963 downto 0);
                        buf_output_r(1002 downto 964) <= data_in(38 downto 0);
                        buf_input_r (24 downto 0)    <= data_in(63 downto 39);
                        bits_in_buffer               <= 25;
                    when 965 =>
                        buf_output_r(964 downto 0)   <= buf_input_r(964 downto 0);
                        buf_output_r(1002 downto 965) <= data_in(37 downto 0);
                        buf_input_r (25 downto 0)    <= data_in(63 downto 38);
                        bits_in_buffer               <= 26;
                    when 966 =>
                        buf_output_r(965 downto 0)   <= buf_input_r(965 downto 0);
                        buf_output_r(1002 downto 966) <= data_in(36 downto 0);
                        buf_input_r (26 downto 0)    <= data_in(63 downto 37);
                        bits_in_buffer               <= 27;
                    when 967 =>
                        buf_output_r(966 downto 0)   <= buf_input_r(966 downto 0);
                        buf_output_r(1002 downto 967) <= data_in(35 downto 0);
                        buf_input_r (27 downto 0)    <= data_in(63 downto 36);
                        bits_in_buffer               <= 28;
                    when 968 =>
                        buf_output_r(967 downto 0)   <= buf_input_r(967 downto 0);
                        buf_output_r(1002 downto 968) <= data_in(34 downto 0);
                        buf_input_r (28 downto 0)    <= data_in(63 downto 35);
                        bits_in_buffer               <= 29;
                    when 969 =>
                        buf_output_r(968 downto 0)   <= buf_input_r(968 downto 0);
                        buf_output_r(1002 downto 969) <= data_in(33 downto 0);
                        buf_input_r (29 downto 0)    <= data_in(63 downto 34);
                        bits_in_buffer               <= 30;
                    when 970 =>
                        buf_output_r(969 downto 0)   <= buf_input_r(969 downto 0);
                        buf_output_r(1002 downto 970) <= data_in(32 downto 0);
                        buf_input_r (30 downto 0)    <= data_in(63 downto 33);
                        bits_in_buffer               <= 31;
                    when 971 =>
                        buf_output_r(970 downto 0)   <= buf_input_r(970 downto 0);
                        buf_output_r(1002 downto 971) <= data_in(31 downto 0);
                        buf_input_r (31 downto 0)    <= data_in(63 downto 32);
                        bits_in_buffer               <= 32;
                    when 972 =>
                        buf_output_r(971 downto 0)   <= buf_input_r(971 downto 0);
                        buf_output_r(1002 downto 972) <= data_in(30 downto 0);
                        buf_input_r (32 downto 0)    <= data_in(63 downto 31);
                        bits_in_buffer               <= 33;
                    when 973 =>
                        buf_output_r(972 downto 0)   <= buf_input_r(972 downto 0);
                        buf_output_r(1002 downto 973) <= data_in(29 downto 0);
                        buf_input_r (33 downto 0)    <= data_in(63 downto 30);
                        bits_in_buffer               <= 34;
                    when 974 =>
                        buf_output_r(973 downto 0)   <= buf_input_r(973 downto 0);
                        buf_output_r(1002 downto 974) <= data_in(28 downto 0);
                        buf_input_r (34 downto 0)    <= data_in(63 downto 29);
                        bits_in_buffer               <= 35;
                    when 975 =>
                        buf_output_r(974 downto 0)   <= buf_input_r(974 downto 0);
                        buf_output_r(1002 downto 975) <= data_in(27 downto 0);
                        buf_input_r (35 downto 0)    <= data_in(63 downto 28);
                        bits_in_buffer               <= 36;
                    when 976 =>
                        buf_output_r(975 downto 0)   <= buf_input_r(975 downto 0);
                        buf_output_r(1002 downto 976) <= data_in(26 downto 0);
                        buf_input_r (36 downto 0)    <= data_in(63 downto 27);
                        bits_in_buffer               <= 37;
                    when 977 =>
                        buf_output_r(976 downto 0)   <= buf_input_r(976 downto 0);
                        buf_output_r(1002 downto 977) <= data_in(25 downto 0);
                        buf_input_r (37 downto 0)    <= data_in(63 downto 26);
                        bits_in_buffer               <= 38;
                    when 978 =>
                        buf_output_r(977 downto 0)   <= buf_input_r(977 downto 0);
                        buf_output_r(1002 downto 978) <= data_in(24 downto 0);
                        buf_input_r (38 downto 0)    <= data_in(63 downto 25);
                        bits_in_buffer               <= 39;
                    when 979 =>
                        buf_output_r(978 downto 0)   <= buf_input_r(978 downto 0);
                        buf_output_r(1002 downto 979) <= data_in(23 downto 0);
                        buf_input_r (39 downto 0)    <= data_in(63 downto 24);
                        bits_in_buffer               <= 40;
                    when 980 =>
                        buf_output_r(979 downto 0)   <= buf_input_r(979 downto 0);
                        buf_output_r(1002 downto 980) <= data_in(22 downto 0);
                        buf_input_r (40 downto 0)    <= data_in(63 downto 23);
                        bits_in_buffer               <= 41;
                    when 981 =>
                        buf_output_r(980 downto 0)   <= buf_input_r(980 downto 0);
                        buf_output_r(1002 downto 981) <= data_in(21 downto 0);
                        buf_input_r (41 downto 0)    <= data_in(63 downto 22);
                        bits_in_buffer               <= 42;
                    when 982 =>
                        buf_output_r(981 downto 0)   <= buf_input_r(981 downto 0);
                        buf_output_r(1002 downto 982) <= data_in(20 downto 0);
                        buf_input_r (42 downto 0)    <= data_in(63 downto 21);
                        bits_in_buffer               <= 43;
                    when 983 =>
                        buf_output_r(982 downto 0)   <= buf_input_r(982 downto 0);
                        buf_output_r(1002 downto 983) <= data_in(19 downto 0);
                        buf_input_r (43 downto 0)    <= data_in(63 downto 20);
                        bits_in_buffer               <= 44;
                    when 984 =>
                        buf_output_r(983 downto 0)   <= buf_input_r(983 downto 0);
                        buf_output_r(1002 downto 984) <= data_in(18 downto 0);
                        buf_input_r (44 downto 0)    <= data_in(63 downto 19);
                        bits_in_buffer               <= 45;
                    when 985 =>
                        buf_output_r(984 downto 0)   <= buf_input_r(984 downto 0);
                        buf_output_r(1002 downto 985) <= data_in(17 downto 0);
                        buf_input_r (45 downto 0)    <= data_in(63 downto 18);
                        bits_in_buffer               <= 46;
                    when 986 =>
                        buf_output_r(985 downto 0)   <= buf_input_r(985 downto 0);
                        buf_output_r(1002 downto 986) <= data_in(16 downto 0);
                        buf_input_r (46 downto 0)    <= data_in(63 downto 17);
                        bits_in_buffer               <= 47;
                    when 987 =>
                        buf_output_r(986 downto 0)   <= buf_input_r(986 downto 0);
                        buf_output_r(1002 downto 987) <= data_in(15 downto 0);
                        buf_input_r (47 downto 0)    <= data_in(63 downto 16);
                        bits_in_buffer               <= 48;
                    when 988 =>
                        buf_output_r(987 downto 0)   <= buf_input_r(987 downto 0);
                        buf_output_r(1002 downto 988) <= data_in(14 downto 0);
                        buf_input_r (48 downto 0)    <= data_in(63 downto 15);
                        bits_in_buffer               <= 49;
                    when 989 =>
                        buf_output_r(988 downto 0)   <= buf_input_r(988 downto 0);
                        buf_output_r(1002 downto 989) <= data_in(13 downto 0);
                        buf_input_r (49 downto 0)    <= data_in(63 downto 14);
                        bits_in_buffer               <= 50;
                    when 990 =>
                        buf_output_r(989 downto 0)   <= buf_input_r(989 downto 0);
                        buf_output_r(1002 downto 990) <= data_in(12 downto 0);
                        buf_input_r (50 downto 0)    <= data_in(63 downto 13);
                        bits_in_buffer               <= 51;
                    when 991 =>
                        buf_output_r(990 downto 0)   <= buf_input_r(990 downto 0);
                        buf_output_r(1002 downto 991) <= data_in(11 downto 0);
                        buf_input_r (51 downto 0)    <= data_in(63 downto 12);
                        bits_in_buffer               <= 52;
                    when 992 =>
                        buf_output_r(991 downto 0)   <= buf_input_r(991 downto 0);
                        buf_output_r(1002 downto 992) <= data_in(10 downto 0);
                        buf_input_r (52 downto 0)    <= data_in(63 downto 11);
                        bits_in_buffer               <= 53;
                    when 993 =>
                        buf_output_r(992 downto 0)   <= buf_input_r(992 downto 0);
                        buf_output_r(1002 downto 993) <= data_in(9 downto 0);
                        buf_input_r (53 downto 0)    <= data_in(63 downto 10);
                        bits_in_buffer               <= 54;
                    when 994 =>
                        buf_output_r(993 downto 0)   <= buf_input_r(993 downto 0);
                        buf_output_r(1002 downto 994) <= data_in(8 downto 0);
                        buf_input_r (54 downto 0)    <= data_in(63 downto 9);
                        bits_in_buffer               <= 55;
                    when 995 =>
                        buf_output_r(994 downto 0)   <= buf_input_r(994 downto 0);
                        buf_output_r(1002 downto 995) <= data_in(7 downto 0);
                        buf_input_r (55 downto 0)    <= data_in(63 downto 8);
                        bits_in_buffer               <= 56;
                    when 996 =>
                        buf_output_r(995 downto 0)   <= buf_input_r(995 downto 0);
                        buf_output_r(1002 downto 996) <= data_in(6 downto 0);
                        buf_input_r (56 downto 0)    <= data_in(63 downto 7);
                        bits_in_buffer               <= 57;
                    when 997 =>
                        buf_output_r(996 downto 0)   <= buf_input_r(996 downto 0);
                        buf_output_r(1002 downto 997) <= data_in(5 downto 0);
                        buf_input_r (57 downto 0)    <= data_in(63 downto 6);
                        bits_in_buffer               <= 58;
                    when 998 =>
                        buf_output_r(997 downto 0)   <= buf_input_r(997 downto 0);
                        buf_output_r(1002 downto 998) <= data_in(4 downto 0);
                        buf_input_r (58 downto 0)    <= data_in(63 downto 5);
                        bits_in_buffer               <= 59;
                    when 999 =>
                        buf_output_r(998 downto 0)   <= buf_input_r(998 downto 0);
                        buf_output_r(1002 downto 999) <= data_in(3 downto 0);
                        buf_input_r (59 downto 0)    <= data_in(63 downto 4);
                        bits_in_buffer               <= 60;
                    when 1000 =>
                        buf_output_r(999 downto 0)   <= buf_input_r(999 downto 0);
                        buf_output_r(1002 downto 1000) <= data_in(2 downto 0);
                        buf_input_r (60 downto 0)    <= data_in(63 downto 3);
                        bits_in_buffer               <= 61;
                    when 1001 =>
                        buf_output_r(1000 downto 0)  <= buf_input_r(1000 downto 0);
                        buf_output_r(1002 downto 1001) <= data_in(1 downto 0);
                        buf_input_r (61 downto 0)    <= data_in(63 downto 2);
                        bits_in_buffer               <= 62;
                    when 1002 =>
                        buf_output_r(1001 downto 0)  <= buf_input_r(1001 downto 0);
                        buf_output_r(1002 downto 1002) <= data_in(0 downto 0);
                        buf_input_r (62 downto 0)    <= data_in(63 downto 1);
                        bits_in_buffer               <= 63;
                    when others =>
                end case;
            else
                out_rdy_r <= '0';
                case bits_in_buffer is
                    when 0 =>
                        buf_input_r (63 downto 0)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 64;
                    when 1 =>
                        buf_input_r (64 downto 1)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 65;
                    when 2 =>
                        buf_input_r (65 downto 2)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 66;
                    when 3 =>
                        buf_input_r (66 downto 3)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 67;
                    when 4 =>
                        buf_input_r (67 downto 4)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 68;
                    when 5 =>
                        buf_input_r (68 downto 5)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 69;
                    when 6 =>
                        buf_input_r (69 downto 6)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 70;
                    when 7 =>
                        buf_input_r (70 downto 7)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 71;
                    when 8 =>
                        buf_input_r (71 downto 8)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 72;
                    when 9 =>
                        buf_input_r (72 downto 9)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 73;
                    when 10 =>
                        buf_input_r (73 downto 10)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 74;
                    when 11 =>
                        buf_input_r (74 downto 11)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 75;
                    when 12 =>
                        buf_input_r (75 downto 12)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 76;
                    when 13 =>
                        buf_input_r (76 downto 13)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 77;
                    when 14 =>
                        buf_input_r (77 downto 14)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 78;
                    when 15 =>
                        buf_input_r (78 downto 15)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 79;
                    when 16 =>
                        buf_input_r (79 downto 16)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 80;
                    when 17 =>
                        buf_input_r (80 downto 17)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 81;
                    when 18 =>
                        buf_input_r (81 downto 18)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 82;
                    when 19 =>
                        buf_input_r (82 downto 19)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 83;
                    when 20 =>
                        buf_input_r (83 downto 20)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 84;
                    when 21 =>
                        buf_input_r (84 downto 21)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 85;
                    when 22 =>
                        buf_input_r (85 downto 22)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 86;
                    when 23 =>
                        buf_input_r (86 downto 23)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 87;
                    when 24 =>
                        buf_input_r (87 downto 24)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 88;
                    when 25 =>
                        buf_input_r (88 downto 25)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 89;
                    when 26 =>
                        buf_input_r (89 downto 26)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 90;
                    when 27 =>
                        buf_input_r (90 downto 27)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 91;
                    when 28 =>
                        buf_input_r (91 downto 28)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 92;
                    when 29 =>
                        buf_input_r (92 downto 29)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 93;
                    when 30 =>
                        buf_input_r (93 downto 30)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 94;
                    when 31 =>
                        buf_input_r (94 downto 31)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 95;
                    when 32 =>
                        buf_input_r (95 downto 32)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 96;
                    when 33 =>
                        buf_input_r (96 downto 33)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 97;
                    when 34 =>
                        buf_input_r (97 downto 34)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 98;
                    when 35 =>
                        buf_input_r (98 downto 35)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 99;
                    when 36 =>
                        buf_input_r (99 downto 36)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 100;
                    when 37 =>
                        buf_input_r (100 downto 37)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 101;
                    when 38 =>
                        buf_input_r (101 downto 38)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 102;
                    when 39 =>
                        buf_input_r (102 downto 39)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 103;
                    when 40 =>
                        buf_input_r (103 downto 40)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 104;
                    when 41 =>
                        buf_input_r (104 downto 41)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 105;
                    when 42 =>
                        buf_input_r (105 downto 42)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 106;
                    when 43 =>
                        buf_input_r (106 downto 43)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 107;
                    when 44 =>
                        buf_input_r (107 downto 44)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 108;
                    when 45 =>
                        buf_input_r (108 downto 45)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 109;
                    when 46 =>
                        buf_input_r (109 downto 46)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 110;
                    when 47 =>
                        buf_input_r (110 downto 47)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 111;
                    when 48 =>
                        buf_input_r (111 downto 48)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 112;
                    when 49 =>
                        buf_input_r (112 downto 49)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 113;
                    when 50 =>
                        buf_input_r (113 downto 50)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 114;
                    when 51 =>
                        buf_input_r (114 downto 51)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 115;
                    when 52 =>
                        buf_input_r (115 downto 52)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 116;
                    when 53 =>
                        buf_input_r (116 downto 53)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 117;
                    when 54 =>
                        buf_input_r (117 downto 54)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 118;
                    when 55 =>
                        buf_input_r (118 downto 55)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 119;
                    when 56 =>
                        buf_input_r (119 downto 56)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 120;
                    when 57 =>
                        buf_input_r (120 downto 57)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 121;
                    when 58 =>
                        buf_input_r (121 downto 58)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 122;
                    when 59 =>
                        buf_input_r (122 downto 59)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 123;
                    when 60 =>
                        buf_input_r (123 downto 60)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 124;
                    when 61 =>
                        buf_input_r (124 downto 61)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 125;
                    when 62 =>
                        buf_input_r (125 downto 62)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 126;
                    when 63 =>
                        buf_input_r (126 downto 63)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 127;
                    when 64 =>
                        buf_input_r (127 downto 64)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 128;
                    when 65 =>
                        buf_input_r (128 downto 65)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 129;
                    when 66 =>
                        buf_input_r (129 downto 66)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 130;
                    when 67 =>
                        buf_input_r (130 downto 67)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 131;
                    when 68 =>
                        buf_input_r (131 downto 68)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 132;
                    when 69 =>
                        buf_input_r (132 downto 69)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 133;
                    when 70 =>
                        buf_input_r (133 downto 70)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 134;
                    when 71 =>
                        buf_input_r (134 downto 71)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 135;
                    when 72 =>
                        buf_input_r (135 downto 72)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 136;
                    when 73 =>
                        buf_input_r (136 downto 73)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 137;
                    when 74 =>
                        buf_input_r (137 downto 74)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 138;
                    when 75 =>
                        buf_input_r (138 downto 75)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 139;
                    when 76 =>
                        buf_input_r (139 downto 76)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 140;
                    when 77 =>
                        buf_input_r (140 downto 77)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 141;
                    when 78 =>
                        buf_input_r (141 downto 78)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 142;
                    when 79 =>
                        buf_input_r (142 downto 79)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 143;
                    when 80 =>
                        buf_input_r (143 downto 80)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 144;
                    when 81 =>
                        buf_input_r (144 downto 81)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 145;
                    when 82 =>
                        buf_input_r (145 downto 82)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 146;
                    when 83 =>
                        buf_input_r (146 downto 83)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 147;
                    when 84 =>
                        buf_input_r (147 downto 84)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 148;
                    when 85 =>
                        buf_input_r (148 downto 85)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 149;
                    when 86 =>
                        buf_input_r (149 downto 86)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 150;
                    when 87 =>
                        buf_input_r (150 downto 87)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 151;
                    when 88 =>
                        buf_input_r (151 downto 88)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 152;
                    when 89 =>
                        buf_input_r (152 downto 89)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 153;
                    when 90 =>
                        buf_input_r (153 downto 90)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 154;
                    when 91 =>
                        buf_input_r (154 downto 91)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 155;
                    when 92 =>
                        buf_input_r (155 downto 92)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 156;
                    when 93 =>
                        buf_input_r (156 downto 93)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 157;
                    when 94 =>
                        buf_input_r (157 downto 94)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 158;
                    when 95 =>
                        buf_input_r (158 downto 95)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 159;
                    when 96 =>
                        buf_input_r (159 downto 96)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 160;
                    when 97 =>
                        buf_input_r (160 downto 97)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 161;
                    when 98 =>
                        buf_input_r (161 downto 98)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 162;
                    when 99 =>
                        buf_input_r (162 downto 99)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 163;
                    when 100 =>
                        buf_input_r (163 downto 100) <= data_in(63 downto 0);
                        bits_in_buffer               <= 164;
                    when 101 =>
                        buf_input_r (164 downto 101) <= data_in(63 downto 0);
                        bits_in_buffer               <= 165;
                    when 102 =>
                        buf_input_r (165 downto 102) <= data_in(63 downto 0);
                        bits_in_buffer               <= 166;
                    when 103 =>
                        buf_input_r (166 downto 103) <= data_in(63 downto 0);
                        bits_in_buffer               <= 167;
                    when 104 =>
                        buf_input_r (167 downto 104) <= data_in(63 downto 0);
                        bits_in_buffer               <= 168;
                    when 105 =>
                        buf_input_r (168 downto 105) <= data_in(63 downto 0);
                        bits_in_buffer               <= 169;
                    when 106 =>
                        buf_input_r (169 downto 106) <= data_in(63 downto 0);
                        bits_in_buffer               <= 170;
                    when 107 =>
                        buf_input_r (170 downto 107) <= data_in(63 downto 0);
                        bits_in_buffer               <= 171;
                    when 108 =>
                        buf_input_r (171 downto 108) <= data_in(63 downto 0);
                        bits_in_buffer               <= 172;
                    when 109 =>
                        buf_input_r (172 downto 109) <= data_in(63 downto 0);
                        bits_in_buffer               <= 173;
                    when 110 =>
                        buf_input_r (173 downto 110) <= data_in(63 downto 0);
                        bits_in_buffer               <= 174;
                    when 111 =>
                        buf_input_r (174 downto 111) <= data_in(63 downto 0);
                        bits_in_buffer               <= 175;
                    when 112 =>
                        buf_input_r (175 downto 112) <= data_in(63 downto 0);
                        bits_in_buffer               <= 176;
                    when 113 =>
                        buf_input_r (176 downto 113) <= data_in(63 downto 0);
                        bits_in_buffer               <= 177;
                    when 114 =>
                        buf_input_r (177 downto 114) <= data_in(63 downto 0);
                        bits_in_buffer               <= 178;
                    when 115 =>
                        buf_input_r (178 downto 115) <= data_in(63 downto 0);
                        bits_in_buffer               <= 179;
                    when 116 =>
                        buf_input_r (179 downto 116) <= data_in(63 downto 0);
                        bits_in_buffer               <= 180;
                    when 117 =>
                        buf_input_r (180 downto 117) <= data_in(63 downto 0);
                        bits_in_buffer               <= 181;
                    when 118 =>
                        buf_input_r (181 downto 118) <= data_in(63 downto 0);
                        bits_in_buffer               <= 182;
                    when 119 =>
                        buf_input_r (182 downto 119) <= data_in(63 downto 0);
                        bits_in_buffer               <= 183;
                    when 120 =>
                        buf_input_r (183 downto 120) <= data_in(63 downto 0);
                        bits_in_buffer               <= 184;
                    when 121 =>
                        buf_input_r (184 downto 121) <= data_in(63 downto 0);
                        bits_in_buffer               <= 185;
                    when 122 =>
                        buf_input_r (185 downto 122) <= data_in(63 downto 0);
                        bits_in_buffer               <= 186;
                    when 123 =>
                        buf_input_r (186 downto 123) <= data_in(63 downto 0);
                        bits_in_buffer               <= 187;
                    when 124 =>
                        buf_input_r (187 downto 124) <= data_in(63 downto 0);
                        bits_in_buffer               <= 188;
                    when 125 =>
                        buf_input_r (188 downto 125) <= data_in(63 downto 0);
                        bits_in_buffer               <= 189;
                    when 126 =>
                        buf_input_r (189 downto 126) <= data_in(63 downto 0);
                        bits_in_buffer               <= 190;
                    when 127 =>
                        buf_input_r (190 downto 127) <= data_in(63 downto 0);
                        bits_in_buffer               <= 191;
                    when 128 =>
                        buf_input_r (191 downto 128) <= data_in(63 downto 0);
                        bits_in_buffer               <= 192;
                    when 129 =>
                        buf_input_r (192 downto 129) <= data_in(63 downto 0);
                        bits_in_buffer               <= 193;
                    when 130 =>
                        buf_input_r (193 downto 130) <= data_in(63 downto 0);
                        bits_in_buffer               <= 194;
                    when 131 =>
                        buf_input_r (194 downto 131) <= data_in(63 downto 0);
                        bits_in_buffer               <= 195;
                    when 132 =>
                        buf_input_r (195 downto 132) <= data_in(63 downto 0);
                        bits_in_buffer               <= 196;
                    when 133 =>
                        buf_input_r (196 downto 133) <= data_in(63 downto 0);
                        bits_in_buffer               <= 197;
                    when 134 =>
                        buf_input_r (197 downto 134) <= data_in(63 downto 0);
                        bits_in_buffer               <= 198;
                    when 135 =>
                        buf_input_r (198 downto 135) <= data_in(63 downto 0);
                        bits_in_buffer               <= 199;
                    when 136 =>
                        buf_input_r (199 downto 136) <= data_in(63 downto 0);
                        bits_in_buffer               <= 200;
                    when 137 =>
                        buf_input_r (200 downto 137) <= data_in(63 downto 0);
                        bits_in_buffer               <= 201;
                    when 138 =>
                        buf_input_r (201 downto 138) <= data_in(63 downto 0);
                        bits_in_buffer               <= 202;
                    when 139 =>
                        buf_input_r (202 downto 139) <= data_in(63 downto 0);
                        bits_in_buffer               <= 203;
                    when 140 =>
                        buf_input_r (203 downto 140) <= data_in(63 downto 0);
                        bits_in_buffer               <= 204;
                    when 141 =>
                        buf_input_r (204 downto 141) <= data_in(63 downto 0);
                        bits_in_buffer               <= 205;
                    when 142 =>
                        buf_input_r (205 downto 142) <= data_in(63 downto 0);
                        bits_in_buffer               <= 206;
                    when 143 =>
                        buf_input_r (206 downto 143) <= data_in(63 downto 0);
                        bits_in_buffer               <= 207;
                    when 144 =>
                        buf_input_r (207 downto 144) <= data_in(63 downto 0);
                        bits_in_buffer               <= 208;
                    when 145 =>
                        buf_input_r (208 downto 145) <= data_in(63 downto 0);
                        bits_in_buffer               <= 209;
                    when 146 =>
                        buf_input_r (209 downto 146) <= data_in(63 downto 0);
                        bits_in_buffer               <= 210;
                    when 147 =>
                        buf_input_r (210 downto 147) <= data_in(63 downto 0);
                        bits_in_buffer               <= 211;
                    when 148 =>
                        buf_input_r (211 downto 148) <= data_in(63 downto 0);
                        bits_in_buffer               <= 212;
                    when 149 =>
                        buf_input_r (212 downto 149) <= data_in(63 downto 0);
                        bits_in_buffer               <= 213;
                    when 150 =>
                        buf_input_r (213 downto 150) <= data_in(63 downto 0);
                        bits_in_buffer               <= 214;
                    when 151 =>
                        buf_input_r (214 downto 151) <= data_in(63 downto 0);
                        bits_in_buffer               <= 215;
                    when 152 =>
                        buf_input_r (215 downto 152) <= data_in(63 downto 0);
                        bits_in_buffer               <= 216;
                    when 153 =>
                        buf_input_r (216 downto 153) <= data_in(63 downto 0);
                        bits_in_buffer               <= 217;
                    when 154 =>
                        buf_input_r (217 downto 154) <= data_in(63 downto 0);
                        bits_in_buffer               <= 218;
                    when 155 =>
                        buf_input_r (218 downto 155) <= data_in(63 downto 0);
                        bits_in_buffer               <= 219;
                    when 156 =>
                        buf_input_r (219 downto 156) <= data_in(63 downto 0);
                        bits_in_buffer               <= 220;
                    when 157 =>
                        buf_input_r (220 downto 157) <= data_in(63 downto 0);
                        bits_in_buffer               <= 221;
                    when 158 =>
                        buf_input_r (221 downto 158) <= data_in(63 downto 0);
                        bits_in_buffer               <= 222;
                    when 159 =>
                        buf_input_r (222 downto 159) <= data_in(63 downto 0);
                        bits_in_buffer               <= 223;
                    when 160 =>
                        buf_input_r (223 downto 160) <= data_in(63 downto 0);
                        bits_in_buffer               <= 224;
                    when 161 =>
                        buf_input_r (224 downto 161) <= data_in(63 downto 0);
                        bits_in_buffer               <= 225;
                    when 162 =>
                        buf_input_r (225 downto 162) <= data_in(63 downto 0);
                        bits_in_buffer               <= 226;
                    when 163 =>
                        buf_input_r (226 downto 163) <= data_in(63 downto 0);
                        bits_in_buffer               <= 227;
                    when 164 =>
                        buf_input_r (227 downto 164) <= data_in(63 downto 0);
                        bits_in_buffer               <= 228;
                    when 165 =>
                        buf_input_r (228 downto 165) <= data_in(63 downto 0);
                        bits_in_buffer               <= 229;
                    when 166 =>
                        buf_input_r (229 downto 166) <= data_in(63 downto 0);
                        bits_in_buffer               <= 230;
                    when 167 =>
                        buf_input_r (230 downto 167) <= data_in(63 downto 0);
                        bits_in_buffer               <= 231;
                    when 168 =>
                        buf_input_r (231 downto 168) <= data_in(63 downto 0);
                        bits_in_buffer               <= 232;
                    when 169 =>
                        buf_input_r (232 downto 169) <= data_in(63 downto 0);
                        bits_in_buffer               <= 233;
                    when 170 =>
                        buf_input_r (233 downto 170) <= data_in(63 downto 0);
                        bits_in_buffer               <= 234;
                    when 171 =>
                        buf_input_r (234 downto 171) <= data_in(63 downto 0);
                        bits_in_buffer               <= 235;
                    when 172 =>
                        buf_input_r (235 downto 172) <= data_in(63 downto 0);
                        bits_in_buffer               <= 236;
                    when 173 =>
                        buf_input_r (236 downto 173) <= data_in(63 downto 0);
                        bits_in_buffer               <= 237;
                    when 174 =>
                        buf_input_r (237 downto 174) <= data_in(63 downto 0);
                        bits_in_buffer               <= 238;
                    when 175 =>
                        buf_input_r (238 downto 175) <= data_in(63 downto 0);
                        bits_in_buffer               <= 239;
                    when 176 =>
                        buf_input_r (239 downto 176) <= data_in(63 downto 0);
                        bits_in_buffer               <= 240;
                    when 177 =>
                        buf_input_r (240 downto 177) <= data_in(63 downto 0);
                        bits_in_buffer               <= 241;
                    when 178 =>
                        buf_input_r (241 downto 178) <= data_in(63 downto 0);
                        bits_in_buffer               <= 242;
                    when 179 =>
                        buf_input_r (242 downto 179) <= data_in(63 downto 0);
                        bits_in_buffer               <= 243;
                    when 180 =>
                        buf_input_r (243 downto 180) <= data_in(63 downto 0);
                        bits_in_buffer               <= 244;
                    when 181 =>
                        buf_input_r (244 downto 181) <= data_in(63 downto 0);
                        bits_in_buffer               <= 245;
                    when 182 =>
                        buf_input_r (245 downto 182) <= data_in(63 downto 0);
                        bits_in_buffer               <= 246;
                    when 183 =>
                        buf_input_r (246 downto 183) <= data_in(63 downto 0);
                        bits_in_buffer               <= 247;
                    when 184 =>
                        buf_input_r (247 downto 184) <= data_in(63 downto 0);
                        bits_in_buffer               <= 248;
                    when 185 =>
                        buf_input_r (248 downto 185) <= data_in(63 downto 0);
                        bits_in_buffer               <= 249;
                    when 186 =>
                        buf_input_r (249 downto 186) <= data_in(63 downto 0);
                        bits_in_buffer               <= 250;
                    when 187 =>
                        buf_input_r (250 downto 187) <= data_in(63 downto 0);
                        bits_in_buffer               <= 251;
                    when 188 =>
                        buf_input_r (251 downto 188) <= data_in(63 downto 0);
                        bits_in_buffer               <= 252;
                    when 189 =>
                        buf_input_r (252 downto 189) <= data_in(63 downto 0);
                        bits_in_buffer               <= 253;
                    when 190 =>
                        buf_input_r (253 downto 190) <= data_in(63 downto 0);
                        bits_in_buffer               <= 254;
                    when 191 =>
                        buf_input_r (254 downto 191) <= data_in(63 downto 0);
                        bits_in_buffer               <= 255;
                    when 192 =>
                        buf_input_r (255 downto 192) <= data_in(63 downto 0);
                        bits_in_buffer               <= 256;
                    when 193 =>
                        buf_input_r (256 downto 193) <= data_in(63 downto 0);
                        bits_in_buffer               <= 257;
                    when 194 =>
                        buf_input_r (257 downto 194) <= data_in(63 downto 0);
                        bits_in_buffer               <= 258;
                    when 195 =>
                        buf_input_r (258 downto 195) <= data_in(63 downto 0);
                        bits_in_buffer               <= 259;
                    when 196 =>
                        buf_input_r (259 downto 196) <= data_in(63 downto 0);
                        bits_in_buffer               <= 260;
                    when 197 =>
                        buf_input_r (260 downto 197) <= data_in(63 downto 0);
                        bits_in_buffer               <= 261;
                    when 198 =>
                        buf_input_r (261 downto 198) <= data_in(63 downto 0);
                        bits_in_buffer               <= 262;
                    when 199 =>
                        buf_input_r (262 downto 199) <= data_in(63 downto 0);
                        bits_in_buffer               <= 263;
                    when 200 =>
                        buf_input_r (263 downto 200) <= data_in(63 downto 0);
                        bits_in_buffer               <= 264;
                    when 201 =>
                        buf_input_r (264 downto 201) <= data_in(63 downto 0);
                        bits_in_buffer               <= 265;
                    when 202 =>
                        buf_input_r (265 downto 202) <= data_in(63 downto 0);
                        bits_in_buffer               <= 266;
                    when 203 =>
                        buf_input_r (266 downto 203) <= data_in(63 downto 0);
                        bits_in_buffer               <= 267;
                    when 204 =>
                        buf_input_r (267 downto 204) <= data_in(63 downto 0);
                        bits_in_buffer               <= 268;
                    when 205 =>
                        buf_input_r (268 downto 205) <= data_in(63 downto 0);
                        bits_in_buffer               <= 269;
                    when 206 =>
                        buf_input_r (269 downto 206) <= data_in(63 downto 0);
                        bits_in_buffer               <= 270;
                    when 207 =>
                        buf_input_r (270 downto 207) <= data_in(63 downto 0);
                        bits_in_buffer               <= 271;
                    when 208 =>
                        buf_input_r (271 downto 208) <= data_in(63 downto 0);
                        bits_in_buffer               <= 272;
                    when 209 =>
                        buf_input_r (272 downto 209) <= data_in(63 downto 0);
                        bits_in_buffer               <= 273;
                    when 210 =>
                        buf_input_r (273 downto 210) <= data_in(63 downto 0);
                        bits_in_buffer               <= 274;
                    when 211 =>
                        buf_input_r (274 downto 211) <= data_in(63 downto 0);
                        bits_in_buffer               <= 275;
                    when 212 =>
                        buf_input_r (275 downto 212) <= data_in(63 downto 0);
                        bits_in_buffer               <= 276;
                    when 213 =>
                        buf_input_r (276 downto 213) <= data_in(63 downto 0);
                        bits_in_buffer               <= 277;
                    when 214 =>
                        buf_input_r (277 downto 214) <= data_in(63 downto 0);
                        bits_in_buffer               <= 278;
                    when 215 =>
                        buf_input_r (278 downto 215) <= data_in(63 downto 0);
                        bits_in_buffer               <= 279;
                    when 216 =>
                        buf_input_r (279 downto 216) <= data_in(63 downto 0);
                        bits_in_buffer               <= 280;
                    when 217 =>
                        buf_input_r (280 downto 217) <= data_in(63 downto 0);
                        bits_in_buffer               <= 281;
                    when 218 =>
                        buf_input_r (281 downto 218) <= data_in(63 downto 0);
                        bits_in_buffer               <= 282;
                    when 219 =>
                        buf_input_r (282 downto 219) <= data_in(63 downto 0);
                        bits_in_buffer               <= 283;
                    when 220 =>
                        buf_input_r (283 downto 220) <= data_in(63 downto 0);
                        bits_in_buffer               <= 284;
                    when 221 =>
                        buf_input_r (284 downto 221) <= data_in(63 downto 0);
                        bits_in_buffer               <= 285;
                    when 222 =>
                        buf_input_r (285 downto 222) <= data_in(63 downto 0);
                        bits_in_buffer               <= 286;
                    when 223 =>
                        buf_input_r (286 downto 223) <= data_in(63 downto 0);
                        bits_in_buffer               <= 287;
                    when 224 =>
                        buf_input_r (287 downto 224) <= data_in(63 downto 0);
                        bits_in_buffer               <= 288;
                    when 225 =>
                        buf_input_r (288 downto 225) <= data_in(63 downto 0);
                        bits_in_buffer               <= 289;
                    when 226 =>
                        buf_input_r (289 downto 226) <= data_in(63 downto 0);
                        bits_in_buffer               <= 290;
                    when 227 =>
                        buf_input_r (290 downto 227) <= data_in(63 downto 0);
                        bits_in_buffer               <= 291;
                    when 228 =>
                        buf_input_r (291 downto 228) <= data_in(63 downto 0);
                        bits_in_buffer               <= 292;
                    when 229 =>
                        buf_input_r (292 downto 229) <= data_in(63 downto 0);
                        bits_in_buffer               <= 293;
                    when 230 =>
                        buf_input_r (293 downto 230) <= data_in(63 downto 0);
                        bits_in_buffer               <= 294;
                    when 231 =>
                        buf_input_r (294 downto 231) <= data_in(63 downto 0);
                        bits_in_buffer               <= 295;
                    when 232 =>
                        buf_input_r (295 downto 232) <= data_in(63 downto 0);
                        bits_in_buffer               <= 296;
                    when 233 =>
                        buf_input_r (296 downto 233) <= data_in(63 downto 0);
                        bits_in_buffer               <= 297;
                    when 234 =>
                        buf_input_r (297 downto 234) <= data_in(63 downto 0);
                        bits_in_buffer               <= 298;
                    when 235 =>
                        buf_input_r (298 downto 235) <= data_in(63 downto 0);
                        bits_in_buffer               <= 299;
                    when 236 =>
                        buf_input_r (299 downto 236) <= data_in(63 downto 0);
                        bits_in_buffer               <= 300;
                    when 237 =>
                        buf_input_r (300 downto 237) <= data_in(63 downto 0);
                        bits_in_buffer               <= 301;
                    when 238 =>
                        buf_input_r (301 downto 238) <= data_in(63 downto 0);
                        bits_in_buffer               <= 302;
                    when 239 =>
                        buf_input_r (302 downto 239) <= data_in(63 downto 0);
                        bits_in_buffer               <= 303;
                    when 240 =>
                        buf_input_r (303 downto 240) <= data_in(63 downto 0);
                        bits_in_buffer               <= 304;
                    when 241 =>
                        buf_input_r (304 downto 241) <= data_in(63 downto 0);
                        bits_in_buffer               <= 305;
                    when 242 =>
                        buf_input_r (305 downto 242) <= data_in(63 downto 0);
                        bits_in_buffer               <= 306;
                    when 243 =>
                        buf_input_r (306 downto 243) <= data_in(63 downto 0);
                        bits_in_buffer               <= 307;
                    when 244 =>
                        buf_input_r (307 downto 244) <= data_in(63 downto 0);
                        bits_in_buffer               <= 308;
                    when 245 =>
                        buf_input_r (308 downto 245) <= data_in(63 downto 0);
                        bits_in_buffer               <= 309;
                    when 246 =>
                        buf_input_r (309 downto 246) <= data_in(63 downto 0);
                        bits_in_buffer               <= 310;
                    when 247 =>
                        buf_input_r (310 downto 247) <= data_in(63 downto 0);
                        bits_in_buffer               <= 311;
                    when 248 =>
                        buf_input_r (311 downto 248) <= data_in(63 downto 0);
                        bits_in_buffer               <= 312;
                    when 249 =>
                        buf_input_r (312 downto 249) <= data_in(63 downto 0);
                        bits_in_buffer               <= 313;
                    when 250 =>
                        buf_input_r (313 downto 250) <= data_in(63 downto 0);
                        bits_in_buffer               <= 314;
                    when 251 =>
                        buf_input_r (314 downto 251) <= data_in(63 downto 0);
                        bits_in_buffer               <= 315;
                    when 252 =>
                        buf_input_r (315 downto 252) <= data_in(63 downto 0);
                        bits_in_buffer               <= 316;
                    when 253 =>
                        buf_input_r (316 downto 253) <= data_in(63 downto 0);
                        bits_in_buffer               <= 317;
                    when 254 =>
                        buf_input_r (317 downto 254) <= data_in(63 downto 0);
                        bits_in_buffer               <= 318;
                    when 255 =>
                        buf_input_r (318 downto 255) <= data_in(63 downto 0);
                        bits_in_buffer               <= 319;
                    when 256 =>
                        buf_input_r (319 downto 256) <= data_in(63 downto 0);
                        bits_in_buffer               <= 320;
                    when 257 =>
                        buf_input_r (320 downto 257) <= data_in(63 downto 0);
                        bits_in_buffer               <= 321;
                    when 258 =>
                        buf_input_r (321 downto 258) <= data_in(63 downto 0);
                        bits_in_buffer               <= 322;
                    when 259 =>
                        buf_input_r (322 downto 259) <= data_in(63 downto 0);
                        bits_in_buffer               <= 323;
                    when 260 =>
                        buf_input_r (323 downto 260) <= data_in(63 downto 0);
                        bits_in_buffer               <= 324;
                    when 261 =>
                        buf_input_r (324 downto 261) <= data_in(63 downto 0);
                        bits_in_buffer               <= 325;
                    when 262 =>
                        buf_input_r (325 downto 262) <= data_in(63 downto 0);
                        bits_in_buffer               <= 326;
                    when 263 =>
                        buf_input_r (326 downto 263) <= data_in(63 downto 0);
                        bits_in_buffer               <= 327;
                    when 264 =>
                        buf_input_r (327 downto 264) <= data_in(63 downto 0);
                        bits_in_buffer               <= 328;
                    when 265 =>
                        buf_input_r (328 downto 265) <= data_in(63 downto 0);
                        bits_in_buffer               <= 329;
                    when 266 =>
                        buf_input_r (329 downto 266) <= data_in(63 downto 0);
                        bits_in_buffer               <= 330;
                    when 267 =>
                        buf_input_r (330 downto 267) <= data_in(63 downto 0);
                        bits_in_buffer               <= 331;
                    when 268 =>
                        buf_input_r (331 downto 268) <= data_in(63 downto 0);
                        bits_in_buffer               <= 332;
                    when 269 =>
                        buf_input_r (332 downto 269) <= data_in(63 downto 0);
                        bits_in_buffer               <= 333;
                    when 270 =>
                        buf_input_r (333 downto 270) <= data_in(63 downto 0);
                        bits_in_buffer               <= 334;
                    when 271 =>
                        buf_input_r (334 downto 271) <= data_in(63 downto 0);
                        bits_in_buffer               <= 335;
                    when 272 =>
                        buf_input_r (335 downto 272) <= data_in(63 downto 0);
                        bits_in_buffer               <= 336;
                    when 273 =>
                        buf_input_r (336 downto 273) <= data_in(63 downto 0);
                        bits_in_buffer               <= 337;
                    when 274 =>
                        buf_input_r (337 downto 274) <= data_in(63 downto 0);
                        bits_in_buffer               <= 338;
                    when 275 =>
                        buf_input_r (338 downto 275) <= data_in(63 downto 0);
                        bits_in_buffer               <= 339;
                    when 276 =>
                        buf_input_r (339 downto 276) <= data_in(63 downto 0);
                        bits_in_buffer               <= 340;
                    when 277 =>
                        buf_input_r (340 downto 277) <= data_in(63 downto 0);
                        bits_in_buffer               <= 341;
                    when 278 =>
                        buf_input_r (341 downto 278) <= data_in(63 downto 0);
                        bits_in_buffer               <= 342;
                    when 279 =>
                        buf_input_r (342 downto 279) <= data_in(63 downto 0);
                        bits_in_buffer               <= 343;
                    when 280 =>
                        buf_input_r (343 downto 280) <= data_in(63 downto 0);
                        bits_in_buffer               <= 344;
                    when 281 =>
                        buf_input_r (344 downto 281) <= data_in(63 downto 0);
                        bits_in_buffer               <= 345;
                    when 282 =>
                        buf_input_r (345 downto 282) <= data_in(63 downto 0);
                        bits_in_buffer               <= 346;
                    when 283 =>
                        buf_input_r (346 downto 283) <= data_in(63 downto 0);
                        bits_in_buffer               <= 347;
                    when 284 =>
                        buf_input_r (347 downto 284) <= data_in(63 downto 0);
                        bits_in_buffer               <= 348;
                    when 285 =>
                        buf_input_r (348 downto 285) <= data_in(63 downto 0);
                        bits_in_buffer               <= 349;
                    when 286 =>
                        buf_input_r (349 downto 286) <= data_in(63 downto 0);
                        bits_in_buffer               <= 350;
                    when 287 =>
                        buf_input_r (350 downto 287) <= data_in(63 downto 0);
                        bits_in_buffer               <= 351;
                    when 288 =>
                        buf_input_r (351 downto 288) <= data_in(63 downto 0);
                        bits_in_buffer               <= 352;
                    when 289 =>
                        buf_input_r (352 downto 289) <= data_in(63 downto 0);
                        bits_in_buffer               <= 353;
                    when 290 =>
                        buf_input_r (353 downto 290) <= data_in(63 downto 0);
                        bits_in_buffer               <= 354;
                    when 291 =>
                        buf_input_r (354 downto 291) <= data_in(63 downto 0);
                        bits_in_buffer               <= 355;
                    when 292 =>
                        buf_input_r (355 downto 292) <= data_in(63 downto 0);
                        bits_in_buffer               <= 356;
                    when 293 =>
                        buf_input_r (356 downto 293) <= data_in(63 downto 0);
                        bits_in_buffer               <= 357;
                    when 294 =>
                        buf_input_r (357 downto 294) <= data_in(63 downto 0);
                        bits_in_buffer               <= 358;
                    when 295 =>
                        buf_input_r (358 downto 295) <= data_in(63 downto 0);
                        bits_in_buffer               <= 359;
                    when 296 =>
                        buf_input_r (359 downto 296) <= data_in(63 downto 0);
                        bits_in_buffer               <= 360;
                    when 297 =>
                        buf_input_r (360 downto 297) <= data_in(63 downto 0);
                        bits_in_buffer               <= 361;
                    when 298 =>
                        buf_input_r (361 downto 298) <= data_in(63 downto 0);
                        bits_in_buffer               <= 362;
                    when 299 =>
                        buf_input_r (362 downto 299) <= data_in(63 downto 0);
                        bits_in_buffer               <= 363;
                    when 300 =>
                        buf_input_r (363 downto 300) <= data_in(63 downto 0);
                        bits_in_buffer               <= 364;
                    when 301 =>
                        buf_input_r (364 downto 301) <= data_in(63 downto 0);
                        bits_in_buffer               <= 365;
                    when 302 =>
                        buf_input_r (365 downto 302) <= data_in(63 downto 0);
                        bits_in_buffer               <= 366;
                    when 303 =>
                        buf_input_r (366 downto 303) <= data_in(63 downto 0);
                        bits_in_buffer               <= 367;
                    when 304 =>
                        buf_input_r (367 downto 304) <= data_in(63 downto 0);
                        bits_in_buffer               <= 368;
                    when 305 =>
                        buf_input_r (368 downto 305) <= data_in(63 downto 0);
                        bits_in_buffer               <= 369;
                    when 306 =>
                        buf_input_r (369 downto 306) <= data_in(63 downto 0);
                        bits_in_buffer               <= 370;
                    when 307 =>
                        buf_input_r (370 downto 307) <= data_in(63 downto 0);
                        bits_in_buffer               <= 371;
                    when 308 =>
                        buf_input_r (371 downto 308) <= data_in(63 downto 0);
                        bits_in_buffer               <= 372;
                    when 309 =>
                        buf_input_r (372 downto 309) <= data_in(63 downto 0);
                        bits_in_buffer               <= 373;
                    when 310 =>
                        buf_input_r (373 downto 310) <= data_in(63 downto 0);
                        bits_in_buffer               <= 374;
                    when 311 =>
                        buf_input_r (374 downto 311) <= data_in(63 downto 0);
                        bits_in_buffer               <= 375;
                    when 312 =>
                        buf_input_r (375 downto 312) <= data_in(63 downto 0);
                        bits_in_buffer               <= 376;
                    when 313 =>
                        buf_input_r (376 downto 313) <= data_in(63 downto 0);
                        bits_in_buffer               <= 377;
                    when 314 =>
                        buf_input_r (377 downto 314) <= data_in(63 downto 0);
                        bits_in_buffer               <= 378;
                    when 315 =>
                        buf_input_r (378 downto 315) <= data_in(63 downto 0);
                        bits_in_buffer               <= 379;
                    when 316 =>
                        buf_input_r (379 downto 316) <= data_in(63 downto 0);
                        bits_in_buffer               <= 380;
                    when 317 =>
                        buf_input_r (380 downto 317) <= data_in(63 downto 0);
                        bits_in_buffer               <= 381;
                    when 318 =>
                        buf_input_r (381 downto 318) <= data_in(63 downto 0);
                        bits_in_buffer               <= 382;
                    when 319 =>
                        buf_input_r (382 downto 319) <= data_in(63 downto 0);
                        bits_in_buffer               <= 383;
                    when 320 =>
                        buf_input_r (383 downto 320) <= data_in(63 downto 0);
                        bits_in_buffer               <= 384;
                    when 321 =>
                        buf_input_r (384 downto 321) <= data_in(63 downto 0);
                        bits_in_buffer               <= 385;
                    when 322 =>
                        buf_input_r (385 downto 322) <= data_in(63 downto 0);
                        bits_in_buffer               <= 386;
                    when 323 =>
                        buf_input_r (386 downto 323) <= data_in(63 downto 0);
                        bits_in_buffer               <= 387;
                    when 324 =>
                        buf_input_r (387 downto 324) <= data_in(63 downto 0);
                        bits_in_buffer               <= 388;
                    when 325 =>
                        buf_input_r (388 downto 325) <= data_in(63 downto 0);
                        bits_in_buffer               <= 389;
                    when 326 =>
                        buf_input_r (389 downto 326) <= data_in(63 downto 0);
                        bits_in_buffer               <= 390;
                    when 327 =>
                        buf_input_r (390 downto 327) <= data_in(63 downto 0);
                        bits_in_buffer               <= 391;
                    when 328 =>
                        buf_input_r (391 downto 328) <= data_in(63 downto 0);
                        bits_in_buffer               <= 392;
                    when 329 =>
                        buf_input_r (392 downto 329) <= data_in(63 downto 0);
                        bits_in_buffer               <= 393;
                    when 330 =>
                        buf_input_r (393 downto 330) <= data_in(63 downto 0);
                        bits_in_buffer               <= 394;
                    when 331 =>
                        buf_input_r (394 downto 331) <= data_in(63 downto 0);
                        bits_in_buffer               <= 395;
                    when 332 =>
                        buf_input_r (395 downto 332) <= data_in(63 downto 0);
                        bits_in_buffer               <= 396;
                    when 333 =>
                        buf_input_r (396 downto 333) <= data_in(63 downto 0);
                        bits_in_buffer               <= 397;
                    when 334 =>
                        buf_input_r (397 downto 334) <= data_in(63 downto 0);
                        bits_in_buffer               <= 398;
                    when 335 =>
                        buf_input_r (398 downto 335) <= data_in(63 downto 0);
                        bits_in_buffer               <= 399;
                    when 336 =>
                        buf_input_r (399 downto 336) <= data_in(63 downto 0);
                        bits_in_buffer               <= 400;
                    when 337 =>
                        buf_input_r (400 downto 337) <= data_in(63 downto 0);
                        bits_in_buffer               <= 401;
                    when 338 =>
                        buf_input_r (401 downto 338) <= data_in(63 downto 0);
                        bits_in_buffer               <= 402;
                    when 339 =>
                        buf_input_r (402 downto 339) <= data_in(63 downto 0);
                        bits_in_buffer               <= 403;
                    when 340 =>
                        buf_input_r (403 downto 340) <= data_in(63 downto 0);
                        bits_in_buffer               <= 404;
                    when 341 =>
                        buf_input_r (404 downto 341) <= data_in(63 downto 0);
                        bits_in_buffer               <= 405;
                    when 342 =>
                        buf_input_r (405 downto 342) <= data_in(63 downto 0);
                        bits_in_buffer               <= 406;
                    when 343 =>
                        buf_input_r (406 downto 343) <= data_in(63 downto 0);
                        bits_in_buffer               <= 407;
                    when 344 =>
                        buf_input_r (407 downto 344) <= data_in(63 downto 0);
                        bits_in_buffer               <= 408;
                    when 345 =>
                        buf_input_r (408 downto 345) <= data_in(63 downto 0);
                        bits_in_buffer               <= 409;
                    when 346 =>
                        buf_input_r (409 downto 346) <= data_in(63 downto 0);
                        bits_in_buffer               <= 410;
                    when 347 =>
                        buf_input_r (410 downto 347) <= data_in(63 downto 0);
                        bits_in_buffer               <= 411;
                    when 348 =>
                        buf_input_r (411 downto 348) <= data_in(63 downto 0);
                        bits_in_buffer               <= 412;
                    when 349 =>
                        buf_input_r (412 downto 349) <= data_in(63 downto 0);
                        bits_in_buffer               <= 413;
                    when 350 =>
                        buf_input_r (413 downto 350) <= data_in(63 downto 0);
                        bits_in_buffer               <= 414;
                    when 351 =>
                        buf_input_r (414 downto 351) <= data_in(63 downto 0);
                        bits_in_buffer               <= 415;
                    when 352 =>
                        buf_input_r (415 downto 352) <= data_in(63 downto 0);
                        bits_in_buffer               <= 416;
                    when 353 =>
                        buf_input_r (416 downto 353) <= data_in(63 downto 0);
                        bits_in_buffer               <= 417;
                    when 354 =>
                        buf_input_r (417 downto 354) <= data_in(63 downto 0);
                        bits_in_buffer               <= 418;
                    when 355 =>
                        buf_input_r (418 downto 355) <= data_in(63 downto 0);
                        bits_in_buffer               <= 419;
                    when 356 =>
                        buf_input_r (419 downto 356) <= data_in(63 downto 0);
                        bits_in_buffer               <= 420;
                    when 357 =>
                        buf_input_r (420 downto 357) <= data_in(63 downto 0);
                        bits_in_buffer               <= 421;
                    when 358 =>
                        buf_input_r (421 downto 358) <= data_in(63 downto 0);
                        bits_in_buffer               <= 422;
                    when 359 =>
                        buf_input_r (422 downto 359) <= data_in(63 downto 0);
                        bits_in_buffer               <= 423;
                    when 360 =>
                        buf_input_r (423 downto 360) <= data_in(63 downto 0);
                        bits_in_buffer               <= 424;
                    when 361 =>
                        buf_input_r (424 downto 361) <= data_in(63 downto 0);
                        bits_in_buffer               <= 425;
                    when 362 =>
                        buf_input_r (425 downto 362) <= data_in(63 downto 0);
                        bits_in_buffer               <= 426;
                    when 363 =>
                        buf_input_r (426 downto 363) <= data_in(63 downto 0);
                        bits_in_buffer               <= 427;
                    when 364 =>
                        buf_input_r (427 downto 364) <= data_in(63 downto 0);
                        bits_in_buffer               <= 428;
                    when 365 =>
                        buf_input_r (428 downto 365) <= data_in(63 downto 0);
                        bits_in_buffer               <= 429;
                    when 366 =>
                        buf_input_r (429 downto 366) <= data_in(63 downto 0);
                        bits_in_buffer               <= 430;
                    when 367 =>
                        buf_input_r (430 downto 367) <= data_in(63 downto 0);
                        bits_in_buffer               <= 431;
                    when 368 =>
                        buf_input_r (431 downto 368) <= data_in(63 downto 0);
                        bits_in_buffer               <= 432;
                    when 369 =>
                        buf_input_r (432 downto 369) <= data_in(63 downto 0);
                        bits_in_buffer               <= 433;
                    when 370 =>
                        buf_input_r (433 downto 370) <= data_in(63 downto 0);
                        bits_in_buffer               <= 434;
                    when 371 =>
                        buf_input_r (434 downto 371) <= data_in(63 downto 0);
                        bits_in_buffer               <= 435;
                    when 372 =>
                        buf_input_r (435 downto 372) <= data_in(63 downto 0);
                        bits_in_buffer               <= 436;
                    when 373 =>
                        buf_input_r (436 downto 373) <= data_in(63 downto 0);
                        bits_in_buffer               <= 437;
                    when 374 =>
                        buf_input_r (437 downto 374) <= data_in(63 downto 0);
                        bits_in_buffer               <= 438;
                    when 375 =>
                        buf_input_r (438 downto 375) <= data_in(63 downto 0);
                        bits_in_buffer               <= 439;
                    when 376 =>
                        buf_input_r (439 downto 376) <= data_in(63 downto 0);
                        bits_in_buffer               <= 440;
                    when 377 =>
                        buf_input_r (440 downto 377) <= data_in(63 downto 0);
                        bits_in_buffer               <= 441;
                    when 378 =>
                        buf_input_r (441 downto 378) <= data_in(63 downto 0);
                        bits_in_buffer               <= 442;
                    when 379 =>
                        buf_input_r (442 downto 379) <= data_in(63 downto 0);
                        bits_in_buffer               <= 443;
                    when 380 =>
                        buf_input_r (443 downto 380) <= data_in(63 downto 0);
                        bits_in_buffer               <= 444;
                    when 381 =>
                        buf_input_r (444 downto 381) <= data_in(63 downto 0);
                        bits_in_buffer               <= 445;
                    when 382 =>
                        buf_input_r (445 downto 382) <= data_in(63 downto 0);
                        bits_in_buffer               <= 446;
                    when 383 =>
                        buf_input_r (446 downto 383) <= data_in(63 downto 0);
                        bits_in_buffer               <= 447;
                    when 384 =>
                        buf_input_r (447 downto 384) <= data_in(63 downto 0);
                        bits_in_buffer               <= 448;
                    when 385 =>
                        buf_input_r (448 downto 385) <= data_in(63 downto 0);
                        bits_in_buffer               <= 449;
                    when 386 =>
                        buf_input_r (449 downto 386) <= data_in(63 downto 0);
                        bits_in_buffer               <= 450;
                    when 387 =>
                        buf_input_r (450 downto 387) <= data_in(63 downto 0);
                        bits_in_buffer               <= 451;
                    when 388 =>
                        buf_input_r (451 downto 388) <= data_in(63 downto 0);
                        bits_in_buffer               <= 452;
                    when 389 =>
                        buf_input_r (452 downto 389) <= data_in(63 downto 0);
                        bits_in_buffer               <= 453;
                    when 390 =>
                        buf_input_r (453 downto 390) <= data_in(63 downto 0);
                        bits_in_buffer               <= 454;
                    when 391 =>
                        buf_input_r (454 downto 391) <= data_in(63 downto 0);
                        bits_in_buffer               <= 455;
                    when 392 =>
                        buf_input_r (455 downto 392) <= data_in(63 downto 0);
                        bits_in_buffer               <= 456;
                    when 393 =>
                        buf_input_r (456 downto 393) <= data_in(63 downto 0);
                        bits_in_buffer               <= 457;
                    when 394 =>
                        buf_input_r (457 downto 394) <= data_in(63 downto 0);
                        bits_in_buffer               <= 458;
                    when 395 =>
                        buf_input_r (458 downto 395) <= data_in(63 downto 0);
                        bits_in_buffer               <= 459;
                    when 396 =>
                        buf_input_r (459 downto 396) <= data_in(63 downto 0);
                        bits_in_buffer               <= 460;
                    when 397 =>
                        buf_input_r (460 downto 397) <= data_in(63 downto 0);
                        bits_in_buffer               <= 461;
                    when 398 =>
                        buf_input_r (461 downto 398) <= data_in(63 downto 0);
                        bits_in_buffer               <= 462;
                    when 399 =>
                        buf_input_r (462 downto 399) <= data_in(63 downto 0);
                        bits_in_buffer               <= 463;
                    when 400 =>
                        buf_input_r (463 downto 400) <= data_in(63 downto 0);
                        bits_in_buffer               <= 464;
                    when 401 =>
                        buf_input_r (464 downto 401) <= data_in(63 downto 0);
                        bits_in_buffer               <= 465;
                    when 402 =>
                        buf_input_r (465 downto 402) <= data_in(63 downto 0);
                        bits_in_buffer               <= 466;
                    when 403 =>
                        buf_input_r (466 downto 403) <= data_in(63 downto 0);
                        bits_in_buffer               <= 467;
                    when 404 =>
                        buf_input_r (467 downto 404) <= data_in(63 downto 0);
                        bits_in_buffer               <= 468;
                    when 405 =>
                        buf_input_r (468 downto 405) <= data_in(63 downto 0);
                        bits_in_buffer               <= 469;
                    when 406 =>
                        buf_input_r (469 downto 406) <= data_in(63 downto 0);
                        bits_in_buffer               <= 470;
                    when 407 =>
                        buf_input_r (470 downto 407) <= data_in(63 downto 0);
                        bits_in_buffer               <= 471;
                    when 408 =>
                        buf_input_r (471 downto 408) <= data_in(63 downto 0);
                        bits_in_buffer               <= 472;
                    when 409 =>
                        buf_input_r (472 downto 409) <= data_in(63 downto 0);
                        bits_in_buffer               <= 473;
                    when 410 =>
                        buf_input_r (473 downto 410) <= data_in(63 downto 0);
                        bits_in_buffer               <= 474;
                    when 411 =>
                        buf_input_r (474 downto 411) <= data_in(63 downto 0);
                        bits_in_buffer               <= 475;
                    when 412 =>
                        buf_input_r (475 downto 412) <= data_in(63 downto 0);
                        bits_in_buffer               <= 476;
                    when 413 =>
                        buf_input_r (476 downto 413) <= data_in(63 downto 0);
                        bits_in_buffer               <= 477;
                    when 414 =>
                        buf_input_r (477 downto 414) <= data_in(63 downto 0);
                        bits_in_buffer               <= 478;
                    when 415 =>
                        buf_input_r (478 downto 415) <= data_in(63 downto 0);
                        bits_in_buffer               <= 479;
                    when 416 =>
                        buf_input_r (479 downto 416) <= data_in(63 downto 0);
                        bits_in_buffer               <= 480;
                    when 417 =>
                        buf_input_r (480 downto 417) <= data_in(63 downto 0);
                        bits_in_buffer               <= 481;
                    when 418 =>
                        buf_input_r (481 downto 418) <= data_in(63 downto 0);
                        bits_in_buffer               <= 482;
                    when 419 =>
                        buf_input_r (482 downto 419) <= data_in(63 downto 0);
                        bits_in_buffer               <= 483;
                    when 420 =>
                        buf_input_r (483 downto 420) <= data_in(63 downto 0);
                        bits_in_buffer               <= 484;
                    when 421 =>
                        buf_input_r (484 downto 421) <= data_in(63 downto 0);
                        bits_in_buffer               <= 485;
                    when 422 =>
                        buf_input_r (485 downto 422) <= data_in(63 downto 0);
                        bits_in_buffer               <= 486;
                    when 423 =>
                        buf_input_r (486 downto 423) <= data_in(63 downto 0);
                        bits_in_buffer               <= 487;
                    when 424 =>
                        buf_input_r (487 downto 424) <= data_in(63 downto 0);
                        bits_in_buffer               <= 488;
                    when 425 =>
                        buf_input_r (488 downto 425) <= data_in(63 downto 0);
                        bits_in_buffer               <= 489;
                    when 426 =>
                        buf_input_r (489 downto 426) <= data_in(63 downto 0);
                        bits_in_buffer               <= 490;
                    when 427 =>
                        buf_input_r (490 downto 427) <= data_in(63 downto 0);
                        bits_in_buffer               <= 491;
                    when 428 =>
                        buf_input_r (491 downto 428) <= data_in(63 downto 0);
                        bits_in_buffer               <= 492;
                    when 429 =>
                        buf_input_r (492 downto 429) <= data_in(63 downto 0);
                        bits_in_buffer               <= 493;
                    when 430 =>
                        buf_input_r (493 downto 430) <= data_in(63 downto 0);
                        bits_in_buffer               <= 494;
                    when 431 =>
                        buf_input_r (494 downto 431) <= data_in(63 downto 0);
                        bits_in_buffer               <= 495;
                    when 432 =>
                        buf_input_r (495 downto 432) <= data_in(63 downto 0);
                        bits_in_buffer               <= 496;
                    when 433 =>
                        buf_input_r (496 downto 433) <= data_in(63 downto 0);
                        bits_in_buffer               <= 497;
                    when 434 =>
                        buf_input_r (497 downto 434) <= data_in(63 downto 0);
                        bits_in_buffer               <= 498;
                    when 435 =>
                        buf_input_r (498 downto 435) <= data_in(63 downto 0);
                        bits_in_buffer               <= 499;
                    when 436 =>
                        buf_input_r (499 downto 436) <= data_in(63 downto 0);
                        bits_in_buffer               <= 500;
                    when 437 =>
                        buf_input_r (500 downto 437) <= data_in(63 downto 0);
                        bits_in_buffer               <= 501;
                    when 438 =>
                        buf_input_r (501 downto 438) <= data_in(63 downto 0);
                        bits_in_buffer               <= 502;
                    when 439 =>
                        buf_input_r (502 downto 439) <= data_in(63 downto 0);
                        bits_in_buffer               <= 503;
                    when 440 =>
                        buf_input_r (503 downto 440) <= data_in(63 downto 0);
                        bits_in_buffer               <= 504;
                    when 441 =>
                        buf_input_r (504 downto 441) <= data_in(63 downto 0);
                        bits_in_buffer               <= 505;
                    when 442 =>
                        buf_input_r (505 downto 442) <= data_in(63 downto 0);
                        bits_in_buffer               <= 506;
                    when 443 =>
                        buf_input_r (506 downto 443) <= data_in(63 downto 0);
                        bits_in_buffer               <= 507;
                    when 444 =>
                        buf_input_r (507 downto 444) <= data_in(63 downto 0);
                        bits_in_buffer               <= 508;
                    when 445 =>
                        buf_input_r (508 downto 445) <= data_in(63 downto 0);
                        bits_in_buffer               <= 509;
                    when 446 =>
                        buf_input_r (509 downto 446) <= data_in(63 downto 0);
                        bits_in_buffer               <= 510;
                    when 447 =>
                        buf_input_r (510 downto 447) <= data_in(63 downto 0);
                        bits_in_buffer               <= 511;
                    when 448 =>
                        buf_input_r (511 downto 448) <= data_in(63 downto 0);
                        bits_in_buffer               <= 512;
                    when 449 =>
                        buf_input_r (512 downto 449) <= data_in(63 downto 0);
                        bits_in_buffer               <= 513;
                    when 450 =>
                        buf_input_r (513 downto 450) <= data_in(63 downto 0);
                        bits_in_buffer               <= 514;
                    when 451 =>
                        buf_input_r (514 downto 451) <= data_in(63 downto 0);
                        bits_in_buffer               <= 515;
                    when 452 =>
                        buf_input_r (515 downto 452) <= data_in(63 downto 0);
                        bits_in_buffer               <= 516;
                    when 453 =>
                        buf_input_r (516 downto 453) <= data_in(63 downto 0);
                        bits_in_buffer               <= 517;
                    when 454 =>
                        buf_input_r (517 downto 454) <= data_in(63 downto 0);
                        bits_in_buffer               <= 518;
                    when 455 =>
                        buf_input_r (518 downto 455) <= data_in(63 downto 0);
                        bits_in_buffer               <= 519;
                    when 456 =>
                        buf_input_r (519 downto 456) <= data_in(63 downto 0);
                        bits_in_buffer               <= 520;
                    when 457 =>
                        buf_input_r (520 downto 457) <= data_in(63 downto 0);
                        bits_in_buffer               <= 521;
                    when 458 =>
                        buf_input_r (521 downto 458) <= data_in(63 downto 0);
                        bits_in_buffer               <= 522;
                    when 459 =>
                        buf_input_r (522 downto 459) <= data_in(63 downto 0);
                        bits_in_buffer               <= 523;
                    when 460 =>
                        buf_input_r (523 downto 460) <= data_in(63 downto 0);
                        bits_in_buffer               <= 524;
                    when 461 =>
                        buf_input_r (524 downto 461) <= data_in(63 downto 0);
                        bits_in_buffer               <= 525;
                    when 462 =>
                        buf_input_r (525 downto 462) <= data_in(63 downto 0);
                        bits_in_buffer               <= 526;
                    when 463 =>
                        buf_input_r (526 downto 463) <= data_in(63 downto 0);
                        bits_in_buffer               <= 527;
                    when 464 =>
                        buf_input_r (527 downto 464) <= data_in(63 downto 0);
                        bits_in_buffer               <= 528;
                    when 465 =>
                        buf_input_r (528 downto 465) <= data_in(63 downto 0);
                        bits_in_buffer               <= 529;
                    when 466 =>
                        buf_input_r (529 downto 466) <= data_in(63 downto 0);
                        bits_in_buffer               <= 530;
                    when 467 =>
                        buf_input_r (530 downto 467) <= data_in(63 downto 0);
                        bits_in_buffer               <= 531;
                    when 468 =>
                        buf_input_r (531 downto 468) <= data_in(63 downto 0);
                        bits_in_buffer               <= 532;
                    when 469 =>
                        buf_input_r (532 downto 469) <= data_in(63 downto 0);
                        bits_in_buffer               <= 533;
                    when 470 =>
                        buf_input_r (533 downto 470) <= data_in(63 downto 0);
                        bits_in_buffer               <= 534;
                    when 471 =>
                        buf_input_r (534 downto 471) <= data_in(63 downto 0);
                        bits_in_buffer               <= 535;
                    when 472 =>
                        buf_input_r (535 downto 472) <= data_in(63 downto 0);
                        bits_in_buffer               <= 536;
                    when 473 =>
                        buf_input_r (536 downto 473) <= data_in(63 downto 0);
                        bits_in_buffer               <= 537;
                    when 474 =>
                        buf_input_r (537 downto 474) <= data_in(63 downto 0);
                        bits_in_buffer               <= 538;
                    when 475 =>
                        buf_input_r (538 downto 475) <= data_in(63 downto 0);
                        bits_in_buffer               <= 539;
                    when 476 =>
                        buf_input_r (539 downto 476) <= data_in(63 downto 0);
                        bits_in_buffer               <= 540;
                    when 477 =>
                        buf_input_r (540 downto 477) <= data_in(63 downto 0);
                        bits_in_buffer               <= 541;
                    when 478 =>
                        buf_input_r (541 downto 478) <= data_in(63 downto 0);
                        bits_in_buffer               <= 542;
                    when 479 =>
                        buf_input_r (542 downto 479) <= data_in(63 downto 0);
                        bits_in_buffer               <= 543;
                    when 480 =>
                        buf_input_r (543 downto 480) <= data_in(63 downto 0);
                        bits_in_buffer               <= 544;
                    when 481 =>
                        buf_input_r (544 downto 481) <= data_in(63 downto 0);
                        bits_in_buffer               <= 545;
                    when 482 =>
                        buf_input_r (545 downto 482) <= data_in(63 downto 0);
                        bits_in_buffer               <= 546;
                    when 483 =>
                        buf_input_r (546 downto 483) <= data_in(63 downto 0);
                        bits_in_buffer               <= 547;
                    when 484 =>
                        buf_input_r (547 downto 484) <= data_in(63 downto 0);
                        bits_in_buffer               <= 548;
                    when 485 =>
                        buf_input_r (548 downto 485) <= data_in(63 downto 0);
                        bits_in_buffer               <= 549;
                    when 486 =>
                        buf_input_r (549 downto 486) <= data_in(63 downto 0);
                        bits_in_buffer               <= 550;
                    when 487 =>
                        buf_input_r (550 downto 487) <= data_in(63 downto 0);
                        bits_in_buffer               <= 551;
                    when 488 =>
                        buf_input_r (551 downto 488) <= data_in(63 downto 0);
                        bits_in_buffer               <= 552;
                    when 489 =>
                        buf_input_r (552 downto 489) <= data_in(63 downto 0);
                        bits_in_buffer               <= 553;
                    when 490 =>
                        buf_input_r (553 downto 490) <= data_in(63 downto 0);
                        bits_in_buffer               <= 554;
                    when 491 =>
                        buf_input_r (554 downto 491) <= data_in(63 downto 0);
                        bits_in_buffer               <= 555;
                    when 492 =>
                        buf_input_r (555 downto 492) <= data_in(63 downto 0);
                        bits_in_buffer               <= 556;
                    when 493 =>
                        buf_input_r (556 downto 493) <= data_in(63 downto 0);
                        bits_in_buffer               <= 557;
                    when 494 =>
                        buf_input_r (557 downto 494) <= data_in(63 downto 0);
                        bits_in_buffer               <= 558;
                    when 495 =>
                        buf_input_r (558 downto 495) <= data_in(63 downto 0);
                        bits_in_buffer               <= 559;
                    when 496 =>
                        buf_input_r (559 downto 496) <= data_in(63 downto 0);
                        bits_in_buffer               <= 560;
                    when 497 =>
                        buf_input_r (560 downto 497) <= data_in(63 downto 0);
                        bits_in_buffer               <= 561;
                    when 498 =>
                        buf_input_r (561 downto 498) <= data_in(63 downto 0);
                        bits_in_buffer               <= 562;
                    when 499 =>
                        buf_input_r (562 downto 499) <= data_in(63 downto 0);
                        bits_in_buffer               <= 563;
                    when 500 =>
                        buf_input_r (563 downto 500) <= data_in(63 downto 0);
                        bits_in_buffer               <= 564;
                    when 501 =>
                        buf_input_r (564 downto 501) <= data_in(63 downto 0);
                        bits_in_buffer               <= 565;
                    when 502 =>
                        buf_input_r (565 downto 502) <= data_in(63 downto 0);
                        bits_in_buffer               <= 566;
                    when 503 =>
                        buf_input_r (566 downto 503) <= data_in(63 downto 0);
                        bits_in_buffer               <= 567;
                    when 504 =>
                        buf_input_r (567 downto 504) <= data_in(63 downto 0);
                        bits_in_buffer               <= 568;
                    when 505 =>
                        buf_input_r (568 downto 505) <= data_in(63 downto 0);
                        bits_in_buffer               <= 569;
                    when 506 =>
                        buf_input_r (569 downto 506) <= data_in(63 downto 0);
                        bits_in_buffer               <= 570;
                    when 507 =>
                        buf_input_r (570 downto 507) <= data_in(63 downto 0);
                        bits_in_buffer               <= 571;
                    when 508 =>
                        buf_input_r (571 downto 508) <= data_in(63 downto 0);
                        bits_in_buffer               <= 572;
                    when 509 =>
                        buf_input_r (572 downto 509) <= data_in(63 downto 0);
                        bits_in_buffer               <= 573;
                    when 510 =>
                        buf_input_r (573 downto 510) <= data_in(63 downto 0);
                        bits_in_buffer               <= 574;
                    when 511 =>
                        buf_input_r (574 downto 511) <= data_in(63 downto 0);
                        bits_in_buffer               <= 575;
                    when 512 =>
                        buf_input_r (575 downto 512) <= data_in(63 downto 0);
                        bits_in_buffer               <= 576;
                    when 513 =>
                        buf_input_r (576 downto 513) <= data_in(63 downto 0);
                        bits_in_buffer               <= 577;
                    when 514 =>
                        buf_input_r (577 downto 514) <= data_in(63 downto 0);
                        bits_in_buffer               <= 578;
                    when 515 =>
                        buf_input_r (578 downto 515) <= data_in(63 downto 0);
                        bits_in_buffer               <= 579;
                    when 516 =>
                        buf_input_r (579 downto 516) <= data_in(63 downto 0);
                        bits_in_buffer               <= 580;
                    when 517 =>
                        buf_input_r (580 downto 517) <= data_in(63 downto 0);
                        bits_in_buffer               <= 581;
                    when 518 =>
                        buf_input_r (581 downto 518) <= data_in(63 downto 0);
                        bits_in_buffer               <= 582;
                    when 519 =>
                        buf_input_r (582 downto 519) <= data_in(63 downto 0);
                        bits_in_buffer               <= 583;
                    when 520 =>
                        buf_input_r (583 downto 520) <= data_in(63 downto 0);
                        bits_in_buffer               <= 584;
                    when 521 =>
                        buf_input_r (584 downto 521) <= data_in(63 downto 0);
                        bits_in_buffer               <= 585;
                    when 522 =>
                        buf_input_r (585 downto 522) <= data_in(63 downto 0);
                        bits_in_buffer               <= 586;
                    when 523 =>
                        buf_input_r (586 downto 523) <= data_in(63 downto 0);
                        bits_in_buffer               <= 587;
                    when 524 =>
                        buf_input_r (587 downto 524) <= data_in(63 downto 0);
                        bits_in_buffer               <= 588;
                    when 525 =>
                        buf_input_r (588 downto 525) <= data_in(63 downto 0);
                        bits_in_buffer               <= 589;
                    when 526 =>
                        buf_input_r (589 downto 526) <= data_in(63 downto 0);
                        bits_in_buffer               <= 590;
                    when 527 =>
                        buf_input_r (590 downto 527) <= data_in(63 downto 0);
                        bits_in_buffer               <= 591;
                    when 528 =>
                        buf_input_r (591 downto 528) <= data_in(63 downto 0);
                        bits_in_buffer               <= 592;
                    when 529 =>
                        buf_input_r (592 downto 529) <= data_in(63 downto 0);
                        bits_in_buffer               <= 593;
                    when 530 =>
                        buf_input_r (593 downto 530) <= data_in(63 downto 0);
                        bits_in_buffer               <= 594;
                    when 531 =>
                        buf_input_r (594 downto 531) <= data_in(63 downto 0);
                        bits_in_buffer               <= 595;
                    when 532 =>
                        buf_input_r (595 downto 532) <= data_in(63 downto 0);
                        bits_in_buffer               <= 596;
                    when 533 =>
                        buf_input_r (596 downto 533) <= data_in(63 downto 0);
                        bits_in_buffer               <= 597;
                    when 534 =>
                        buf_input_r (597 downto 534) <= data_in(63 downto 0);
                        bits_in_buffer               <= 598;
                    when 535 =>
                        buf_input_r (598 downto 535) <= data_in(63 downto 0);
                        bits_in_buffer               <= 599;
                    when 536 =>
                        buf_input_r (599 downto 536) <= data_in(63 downto 0);
                        bits_in_buffer               <= 600;
                    when 537 =>
                        buf_input_r (600 downto 537) <= data_in(63 downto 0);
                        bits_in_buffer               <= 601;
                    when 538 =>
                        buf_input_r (601 downto 538) <= data_in(63 downto 0);
                        bits_in_buffer               <= 602;
                    when 539 =>
                        buf_input_r (602 downto 539) <= data_in(63 downto 0);
                        bits_in_buffer               <= 603;
                    when 540 =>
                        buf_input_r (603 downto 540) <= data_in(63 downto 0);
                        bits_in_buffer               <= 604;
                    when 541 =>
                        buf_input_r (604 downto 541) <= data_in(63 downto 0);
                        bits_in_buffer               <= 605;
                    when 542 =>
                        buf_input_r (605 downto 542) <= data_in(63 downto 0);
                        bits_in_buffer               <= 606;
                    when 543 =>
                        buf_input_r (606 downto 543) <= data_in(63 downto 0);
                        bits_in_buffer               <= 607;
                    when 544 =>
                        buf_input_r (607 downto 544) <= data_in(63 downto 0);
                        bits_in_buffer               <= 608;
                    when 545 =>
                        buf_input_r (608 downto 545) <= data_in(63 downto 0);
                        bits_in_buffer               <= 609;
                    when 546 =>
                        buf_input_r (609 downto 546) <= data_in(63 downto 0);
                        bits_in_buffer               <= 610;
                    when 547 =>
                        buf_input_r (610 downto 547) <= data_in(63 downto 0);
                        bits_in_buffer               <= 611;
                    when 548 =>
                        buf_input_r (611 downto 548) <= data_in(63 downto 0);
                        bits_in_buffer               <= 612;
                    when 549 =>
                        buf_input_r (612 downto 549) <= data_in(63 downto 0);
                        bits_in_buffer               <= 613;
                    when 550 =>
                        buf_input_r (613 downto 550) <= data_in(63 downto 0);
                        bits_in_buffer               <= 614;
                    when 551 =>
                        buf_input_r (614 downto 551) <= data_in(63 downto 0);
                        bits_in_buffer               <= 615;
                    when 552 =>
                        buf_input_r (615 downto 552) <= data_in(63 downto 0);
                        bits_in_buffer               <= 616;
                    when 553 =>
                        buf_input_r (616 downto 553) <= data_in(63 downto 0);
                        bits_in_buffer               <= 617;
                    when 554 =>
                        buf_input_r (617 downto 554) <= data_in(63 downto 0);
                        bits_in_buffer               <= 618;
                    when 555 =>
                        buf_input_r (618 downto 555) <= data_in(63 downto 0);
                        bits_in_buffer               <= 619;
                    when 556 =>
                        buf_input_r (619 downto 556) <= data_in(63 downto 0);
                        bits_in_buffer               <= 620;
                    when 557 =>
                        buf_input_r (620 downto 557) <= data_in(63 downto 0);
                        bits_in_buffer               <= 621;
                    when 558 =>
                        buf_input_r (621 downto 558) <= data_in(63 downto 0);
                        bits_in_buffer               <= 622;
                    when 559 =>
                        buf_input_r (622 downto 559) <= data_in(63 downto 0);
                        bits_in_buffer               <= 623;
                    when 560 =>
                        buf_input_r (623 downto 560) <= data_in(63 downto 0);
                        bits_in_buffer               <= 624;
                    when 561 =>
                        buf_input_r (624 downto 561) <= data_in(63 downto 0);
                        bits_in_buffer               <= 625;
                    when 562 =>
                        buf_input_r (625 downto 562) <= data_in(63 downto 0);
                        bits_in_buffer               <= 626;
                    when 563 =>
                        buf_input_r (626 downto 563) <= data_in(63 downto 0);
                        bits_in_buffer               <= 627;
                    when 564 =>
                        buf_input_r (627 downto 564) <= data_in(63 downto 0);
                        bits_in_buffer               <= 628;
                    when 565 =>
                        buf_input_r (628 downto 565) <= data_in(63 downto 0);
                        bits_in_buffer               <= 629;
                    when 566 =>
                        buf_input_r (629 downto 566) <= data_in(63 downto 0);
                        bits_in_buffer               <= 630;
                    when 567 =>
                        buf_input_r (630 downto 567) <= data_in(63 downto 0);
                        bits_in_buffer               <= 631;
                    when 568 =>
                        buf_input_r (631 downto 568) <= data_in(63 downto 0);
                        bits_in_buffer               <= 632;
                    when 569 =>
                        buf_input_r (632 downto 569) <= data_in(63 downto 0);
                        bits_in_buffer               <= 633;
                    when 570 =>
                        buf_input_r (633 downto 570) <= data_in(63 downto 0);
                        bits_in_buffer               <= 634;
                    when 571 =>
                        buf_input_r (634 downto 571) <= data_in(63 downto 0);
                        bits_in_buffer               <= 635;
                    when 572 =>
                        buf_input_r (635 downto 572) <= data_in(63 downto 0);
                        bits_in_buffer               <= 636;
                    when 573 =>
                        buf_input_r (636 downto 573) <= data_in(63 downto 0);
                        bits_in_buffer               <= 637;
                    when 574 =>
                        buf_input_r (637 downto 574) <= data_in(63 downto 0);
                        bits_in_buffer               <= 638;
                    when 575 =>
                        buf_input_r (638 downto 575) <= data_in(63 downto 0);
                        bits_in_buffer               <= 639;
                    when 576 =>
                        buf_input_r (639 downto 576) <= data_in(63 downto 0);
                        bits_in_buffer               <= 640;
                    when 577 =>
                        buf_input_r (640 downto 577) <= data_in(63 downto 0);
                        bits_in_buffer               <= 641;
                    when 578 =>
                        buf_input_r (641 downto 578) <= data_in(63 downto 0);
                        bits_in_buffer               <= 642;
                    when 579 =>
                        buf_input_r (642 downto 579) <= data_in(63 downto 0);
                        bits_in_buffer               <= 643;
                    when 580 =>
                        buf_input_r (643 downto 580) <= data_in(63 downto 0);
                        bits_in_buffer               <= 644;
                    when 581 =>
                        buf_input_r (644 downto 581) <= data_in(63 downto 0);
                        bits_in_buffer               <= 645;
                    when 582 =>
                        buf_input_r (645 downto 582) <= data_in(63 downto 0);
                        bits_in_buffer               <= 646;
                    when 583 =>
                        buf_input_r (646 downto 583) <= data_in(63 downto 0);
                        bits_in_buffer               <= 647;
                    when 584 =>
                        buf_input_r (647 downto 584) <= data_in(63 downto 0);
                        bits_in_buffer               <= 648;
                    when 585 =>
                        buf_input_r (648 downto 585) <= data_in(63 downto 0);
                        bits_in_buffer               <= 649;
                    when 586 =>
                        buf_input_r (649 downto 586) <= data_in(63 downto 0);
                        bits_in_buffer               <= 650;
                    when 587 =>
                        buf_input_r (650 downto 587) <= data_in(63 downto 0);
                        bits_in_buffer               <= 651;
                    when 588 =>
                        buf_input_r (651 downto 588) <= data_in(63 downto 0);
                        bits_in_buffer               <= 652;
                    when 589 =>
                        buf_input_r (652 downto 589) <= data_in(63 downto 0);
                        bits_in_buffer               <= 653;
                    when 590 =>
                        buf_input_r (653 downto 590) <= data_in(63 downto 0);
                        bits_in_buffer               <= 654;
                    when 591 =>
                        buf_input_r (654 downto 591) <= data_in(63 downto 0);
                        bits_in_buffer               <= 655;
                    when 592 =>
                        buf_input_r (655 downto 592) <= data_in(63 downto 0);
                        bits_in_buffer               <= 656;
                    when 593 =>
                        buf_input_r (656 downto 593) <= data_in(63 downto 0);
                        bits_in_buffer               <= 657;
                    when 594 =>
                        buf_input_r (657 downto 594) <= data_in(63 downto 0);
                        bits_in_buffer               <= 658;
                    when 595 =>
                        buf_input_r (658 downto 595) <= data_in(63 downto 0);
                        bits_in_buffer               <= 659;
                    when 596 =>
                        buf_input_r (659 downto 596) <= data_in(63 downto 0);
                        bits_in_buffer               <= 660;
                    when 597 =>
                        buf_input_r (660 downto 597) <= data_in(63 downto 0);
                        bits_in_buffer               <= 661;
                    when 598 =>
                        buf_input_r (661 downto 598) <= data_in(63 downto 0);
                        bits_in_buffer               <= 662;
                    when 599 =>
                        buf_input_r (662 downto 599) <= data_in(63 downto 0);
                        bits_in_buffer               <= 663;
                    when 600 =>
                        buf_input_r (663 downto 600) <= data_in(63 downto 0);
                        bits_in_buffer               <= 664;
                    when 601 =>
                        buf_input_r (664 downto 601) <= data_in(63 downto 0);
                        bits_in_buffer               <= 665;
                    when 602 =>
                        buf_input_r (665 downto 602) <= data_in(63 downto 0);
                        bits_in_buffer               <= 666;
                    when 603 =>
                        buf_input_r (666 downto 603) <= data_in(63 downto 0);
                        bits_in_buffer               <= 667;
                    when 604 =>
                        buf_input_r (667 downto 604) <= data_in(63 downto 0);
                        bits_in_buffer               <= 668;
                    when 605 =>
                        buf_input_r (668 downto 605) <= data_in(63 downto 0);
                        bits_in_buffer               <= 669;
                    when 606 =>
                        buf_input_r (669 downto 606) <= data_in(63 downto 0);
                        bits_in_buffer               <= 670;
                    when 607 =>
                        buf_input_r (670 downto 607) <= data_in(63 downto 0);
                        bits_in_buffer               <= 671;
                    when 608 =>
                        buf_input_r (671 downto 608) <= data_in(63 downto 0);
                        bits_in_buffer               <= 672;
                    when 609 =>
                        buf_input_r (672 downto 609) <= data_in(63 downto 0);
                        bits_in_buffer               <= 673;
                    when 610 =>
                        buf_input_r (673 downto 610) <= data_in(63 downto 0);
                        bits_in_buffer               <= 674;
                    when 611 =>
                        buf_input_r (674 downto 611) <= data_in(63 downto 0);
                        bits_in_buffer               <= 675;
                    when 612 =>
                        buf_input_r (675 downto 612) <= data_in(63 downto 0);
                        bits_in_buffer               <= 676;
                    when 613 =>
                        buf_input_r (676 downto 613) <= data_in(63 downto 0);
                        bits_in_buffer               <= 677;
                    when 614 =>
                        buf_input_r (677 downto 614) <= data_in(63 downto 0);
                        bits_in_buffer               <= 678;
                    when 615 =>
                        buf_input_r (678 downto 615) <= data_in(63 downto 0);
                        bits_in_buffer               <= 679;
                    when 616 =>
                        buf_input_r (679 downto 616) <= data_in(63 downto 0);
                        bits_in_buffer               <= 680;
                    when 617 =>
                        buf_input_r (680 downto 617) <= data_in(63 downto 0);
                        bits_in_buffer               <= 681;
                    when 618 =>
                        buf_input_r (681 downto 618) <= data_in(63 downto 0);
                        bits_in_buffer               <= 682;
                    when 619 =>
                        buf_input_r (682 downto 619) <= data_in(63 downto 0);
                        bits_in_buffer               <= 683;
                    when 620 =>
                        buf_input_r (683 downto 620) <= data_in(63 downto 0);
                        bits_in_buffer               <= 684;
                    when 621 =>
                        buf_input_r (684 downto 621) <= data_in(63 downto 0);
                        bits_in_buffer               <= 685;
                    when 622 =>
                        buf_input_r (685 downto 622) <= data_in(63 downto 0);
                        bits_in_buffer               <= 686;
                    when 623 =>
                        buf_input_r (686 downto 623) <= data_in(63 downto 0);
                        bits_in_buffer               <= 687;
                    when 624 =>
                        buf_input_r (687 downto 624) <= data_in(63 downto 0);
                        bits_in_buffer               <= 688;
                    when 625 =>
                        buf_input_r (688 downto 625) <= data_in(63 downto 0);
                        bits_in_buffer               <= 689;
                    when 626 =>
                        buf_input_r (689 downto 626) <= data_in(63 downto 0);
                        bits_in_buffer               <= 690;
                    when 627 =>
                        buf_input_r (690 downto 627) <= data_in(63 downto 0);
                        bits_in_buffer               <= 691;
                    when 628 =>
                        buf_input_r (691 downto 628) <= data_in(63 downto 0);
                        bits_in_buffer               <= 692;
                    when 629 =>
                        buf_input_r (692 downto 629) <= data_in(63 downto 0);
                        bits_in_buffer               <= 693;
                    when 630 =>
                        buf_input_r (693 downto 630) <= data_in(63 downto 0);
                        bits_in_buffer               <= 694;
                    when 631 =>
                        buf_input_r (694 downto 631) <= data_in(63 downto 0);
                        bits_in_buffer               <= 695;
                    when 632 =>
                        buf_input_r (695 downto 632) <= data_in(63 downto 0);
                        bits_in_buffer               <= 696;
                    when 633 =>
                        buf_input_r (696 downto 633) <= data_in(63 downto 0);
                        bits_in_buffer               <= 697;
                    when 634 =>
                        buf_input_r (697 downto 634) <= data_in(63 downto 0);
                        bits_in_buffer               <= 698;
                    when 635 =>
                        buf_input_r (698 downto 635) <= data_in(63 downto 0);
                        bits_in_buffer               <= 699;
                    when 636 =>
                        buf_input_r (699 downto 636) <= data_in(63 downto 0);
                        bits_in_buffer               <= 700;
                    when 637 =>
                        buf_input_r (700 downto 637) <= data_in(63 downto 0);
                        bits_in_buffer               <= 701;
                    when 638 =>
                        buf_input_r (701 downto 638) <= data_in(63 downto 0);
                        bits_in_buffer               <= 702;
                    when 639 =>
                        buf_input_r (702 downto 639) <= data_in(63 downto 0);
                        bits_in_buffer               <= 703;
                    when 640 =>
                        buf_input_r (703 downto 640) <= data_in(63 downto 0);
                        bits_in_buffer               <= 704;
                    when 641 =>
                        buf_input_r (704 downto 641) <= data_in(63 downto 0);
                        bits_in_buffer               <= 705;
                    when 642 =>
                        buf_input_r (705 downto 642) <= data_in(63 downto 0);
                        bits_in_buffer               <= 706;
                    when 643 =>
                        buf_input_r (706 downto 643) <= data_in(63 downto 0);
                        bits_in_buffer               <= 707;
                    when 644 =>
                        buf_input_r (707 downto 644) <= data_in(63 downto 0);
                        bits_in_buffer               <= 708;
                    when 645 =>
                        buf_input_r (708 downto 645) <= data_in(63 downto 0);
                        bits_in_buffer               <= 709;
                    when 646 =>
                        buf_input_r (709 downto 646) <= data_in(63 downto 0);
                        bits_in_buffer               <= 710;
                    when 647 =>
                        buf_input_r (710 downto 647) <= data_in(63 downto 0);
                        bits_in_buffer               <= 711;
                    when 648 =>
                        buf_input_r (711 downto 648) <= data_in(63 downto 0);
                        bits_in_buffer               <= 712;
                    when 649 =>
                        buf_input_r (712 downto 649) <= data_in(63 downto 0);
                        bits_in_buffer               <= 713;
                    when 650 =>
                        buf_input_r (713 downto 650) <= data_in(63 downto 0);
                        bits_in_buffer               <= 714;
                    when 651 =>
                        buf_input_r (714 downto 651) <= data_in(63 downto 0);
                        bits_in_buffer               <= 715;
                    when 652 =>
                        buf_input_r (715 downto 652) <= data_in(63 downto 0);
                        bits_in_buffer               <= 716;
                    when 653 =>
                        buf_input_r (716 downto 653) <= data_in(63 downto 0);
                        bits_in_buffer               <= 717;
                    when 654 =>
                        buf_input_r (717 downto 654) <= data_in(63 downto 0);
                        bits_in_buffer               <= 718;
                    when 655 =>
                        buf_input_r (718 downto 655) <= data_in(63 downto 0);
                        bits_in_buffer               <= 719;
                    when 656 =>
                        buf_input_r (719 downto 656) <= data_in(63 downto 0);
                        bits_in_buffer               <= 720;
                    when 657 =>
                        buf_input_r (720 downto 657) <= data_in(63 downto 0);
                        bits_in_buffer               <= 721;
                    when 658 =>
                        buf_input_r (721 downto 658) <= data_in(63 downto 0);
                        bits_in_buffer               <= 722;
                    when 659 =>
                        buf_input_r (722 downto 659) <= data_in(63 downto 0);
                        bits_in_buffer               <= 723;
                    when 660 =>
                        buf_input_r (723 downto 660) <= data_in(63 downto 0);
                        bits_in_buffer               <= 724;
                    when 661 =>
                        buf_input_r (724 downto 661) <= data_in(63 downto 0);
                        bits_in_buffer               <= 725;
                    when 662 =>
                        buf_input_r (725 downto 662) <= data_in(63 downto 0);
                        bits_in_buffer               <= 726;
                    when 663 =>
                        buf_input_r (726 downto 663) <= data_in(63 downto 0);
                        bits_in_buffer               <= 727;
                    when 664 =>
                        buf_input_r (727 downto 664) <= data_in(63 downto 0);
                        bits_in_buffer               <= 728;
                    when 665 =>
                        buf_input_r (728 downto 665) <= data_in(63 downto 0);
                        bits_in_buffer               <= 729;
                    when 666 =>
                        buf_input_r (729 downto 666) <= data_in(63 downto 0);
                        bits_in_buffer               <= 730;
                    when 667 =>
                        buf_input_r (730 downto 667) <= data_in(63 downto 0);
                        bits_in_buffer               <= 731;
                    when 668 =>
                        buf_input_r (731 downto 668) <= data_in(63 downto 0);
                        bits_in_buffer               <= 732;
                    when 669 =>
                        buf_input_r (732 downto 669) <= data_in(63 downto 0);
                        bits_in_buffer               <= 733;
                    when 670 =>
                        buf_input_r (733 downto 670) <= data_in(63 downto 0);
                        bits_in_buffer               <= 734;
                    when 671 =>
                        buf_input_r (734 downto 671) <= data_in(63 downto 0);
                        bits_in_buffer               <= 735;
                    when 672 =>
                        buf_input_r (735 downto 672) <= data_in(63 downto 0);
                        bits_in_buffer               <= 736;
                    when 673 =>
                        buf_input_r (736 downto 673) <= data_in(63 downto 0);
                        bits_in_buffer               <= 737;
                    when 674 =>
                        buf_input_r (737 downto 674) <= data_in(63 downto 0);
                        bits_in_buffer               <= 738;
                    when 675 =>
                        buf_input_r (738 downto 675) <= data_in(63 downto 0);
                        bits_in_buffer               <= 739;
                    when 676 =>
                        buf_input_r (739 downto 676) <= data_in(63 downto 0);
                        bits_in_buffer               <= 740;
                    when 677 =>
                        buf_input_r (740 downto 677) <= data_in(63 downto 0);
                        bits_in_buffer               <= 741;
                    when 678 =>
                        buf_input_r (741 downto 678) <= data_in(63 downto 0);
                        bits_in_buffer               <= 742;
                    when 679 =>
                        buf_input_r (742 downto 679) <= data_in(63 downto 0);
                        bits_in_buffer               <= 743;
                    when 680 =>
                        buf_input_r (743 downto 680) <= data_in(63 downto 0);
                        bits_in_buffer               <= 744;
                    when 681 =>
                        buf_input_r (744 downto 681) <= data_in(63 downto 0);
                        bits_in_buffer               <= 745;
                    when 682 =>
                        buf_input_r (745 downto 682) <= data_in(63 downto 0);
                        bits_in_buffer               <= 746;
                    when 683 =>
                        buf_input_r (746 downto 683) <= data_in(63 downto 0);
                        bits_in_buffer               <= 747;
                    when 684 =>
                        buf_input_r (747 downto 684) <= data_in(63 downto 0);
                        bits_in_buffer               <= 748;
                    when 685 =>
                        buf_input_r (748 downto 685) <= data_in(63 downto 0);
                        bits_in_buffer               <= 749;
                    when 686 =>
                        buf_input_r (749 downto 686) <= data_in(63 downto 0);
                        bits_in_buffer               <= 750;
                    when 687 =>
                        buf_input_r (750 downto 687) <= data_in(63 downto 0);
                        bits_in_buffer               <= 751;
                    when 688 =>
                        buf_input_r (751 downto 688) <= data_in(63 downto 0);
                        bits_in_buffer               <= 752;
                    when 689 =>
                        buf_input_r (752 downto 689) <= data_in(63 downto 0);
                        bits_in_buffer               <= 753;
                    when 690 =>
                        buf_input_r (753 downto 690) <= data_in(63 downto 0);
                        bits_in_buffer               <= 754;
                    when 691 =>
                        buf_input_r (754 downto 691) <= data_in(63 downto 0);
                        bits_in_buffer               <= 755;
                    when 692 =>
                        buf_input_r (755 downto 692) <= data_in(63 downto 0);
                        bits_in_buffer               <= 756;
                    when 693 =>
                        buf_input_r (756 downto 693) <= data_in(63 downto 0);
                        bits_in_buffer               <= 757;
                    when 694 =>
                        buf_input_r (757 downto 694) <= data_in(63 downto 0);
                        bits_in_buffer               <= 758;
                    when 695 =>
                        buf_input_r (758 downto 695) <= data_in(63 downto 0);
                        bits_in_buffer               <= 759;
                    when 696 =>
                        buf_input_r (759 downto 696) <= data_in(63 downto 0);
                        bits_in_buffer               <= 760;
                    when 697 =>
                        buf_input_r (760 downto 697) <= data_in(63 downto 0);
                        bits_in_buffer               <= 761;
                    when 698 =>
                        buf_input_r (761 downto 698) <= data_in(63 downto 0);
                        bits_in_buffer               <= 762;
                    when 699 =>
                        buf_input_r (762 downto 699) <= data_in(63 downto 0);
                        bits_in_buffer               <= 763;
                    when 700 =>
                        buf_input_r (763 downto 700) <= data_in(63 downto 0);
                        bits_in_buffer               <= 764;
                    when 701 =>
                        buf_input_r (764 downto 701) <= data_in(63 downto 0);
                        bits_in_buffer               <= 765;
                    when 702 =>
                        buf_input_r (765 downto 702) <= data_in(63 downto 0);
                        bits_in_buffer               <= 766;
                    when 703 =>
                        buf_input_r (766 downto 703) <= data_in(63 downto 0);
                        bits_in_buffer               <= 767;
                    when 704 =>
                        buf_input_r (767 downto 704) <= data_in(63 downto 0);
                        bits_in_buffer               <= 768;
                    when 705 =>
                        buf_input_r (768 downto 705) <= data_in(63 downto 0);
                        bits_in_buffer               <= 769;
                    when 706 =>
                        buf_input_r (769 downto 706) <= data_in(63 downto 0);
                        bits_in_buffer               <= 770;
                    when 707 =>
                        buf_input_r (770 downto 707) <= data_in(63 downto 0);
                        bits_in_buffer               <= 771;
                    when 708 =>
                        buf_input_r (771 downto 708) <= data_in(63 downto 0);
                        bits_in_buffer               <= 772;
                    when 709 =>
                        buf_input_r (772 downto 709) <= data_in(63 downto 0);
                        bits_in_buffer               <= 773;
                    when 710 =>
                        buf_input_r (773 downto 710) <= data_in(63 downto 0);
                        bits_in_buffer               <= 774;
                    when 711 =>
                        buf_input_r (774 downto 711) <= data_in(63 downto 0);
                        bits_in_buffer               <= 775;
                    when 712 =>
                        buf_input_r (775 downto 712) <= data_in(63 downto 0);
                        bits_in_buffer               <= 776;
                    when 713 =>
                        buf_input_r (776 downto 713) <= data_in(63 downto 0);
                        bits_in_buffer               <= 777;
                    when 714 =>
                        buf_input_r (777 downto 714) <= data_in(63 downto 0);
                        bits_in_buffer               <= 778;
                    when 715 =>
                        buf_input_r (778 downto 715) <= data_in(63 downto 0);
                        bits_in_buffer               <= 779;
                    when 716 =>
                        buf_input_r (779 downto 716) <= data_in(63 downto 0);
                        bits_in_buffer               <= 780;
                    when 717 =>
                        buf_input_r (780 downto 717) <= data_in(63 downto 0);
                        bits_in_buffer               <= 781;
                    when 718 =>
                        buf_input_r (781 downto 718) <= data_in(63 downto 0);
                        bits_in_buffer               <= 782;
                    when 719 =>
                        buf_input_r (782 downto 719) <= data_in(63 downto 0);
                        bits_in_buffer               <= 783;
                    when 720 =>
                        buf_input_r (783 downto 720) <= data_in(63 downto 0);
                        bits_in_buffer               <= 784;
                    when 721 =>
                        buf_input_r (784 downto 721) <= data_in(63 downto 0);
                        bits_in_buffer               <= 785;
                    when 722 =>
                        buf_input_r (785 downto 722) <= data_in(63 downto 0);
                        bits_in_buffer               <= 786;
                    when 723 =>
                        buf_input_r (786 downto 723) <= data_in(63 downto 0);
                        bits_in_buffer               <= 787;
                    when 724 =>
                        buf_input_r (787 downto 724) <= data_in(63 downto 0);
                        bits_in_buffer               <= 788;
                    when 725 =>
                        buf_input_r (788 downto 725) <= data_in(63 downto 0);
                        bits_in_buffer               <= 789;
                    when 726 =>
                        buf_input_r (789 downto 726) <= data_in(63 downto 0);
                        bits_in_buffer               <= 790;
                    when 727 =>
                        buf_input_r (790 downto 727) <= data_in(63 downto 0);
                        bits_in_buffer               <= 791;
                    when 728 =>
                        buf_input_r (791 downto 728) <= data_in(63 downto 0);
                        bits_in_buffer               <= 792;
                    when 729 =>
                        buf_input_r (792 downto 729) <= data_in(63 downto 0);
                        bits_in_buffer               <= 793;
                    when 730 =>
                        buf_input_r (793 downto 730) <= data_in(63 downto 0);
                        bits_in_buffer               <= 794;
                    when 731 =>
                        buf_input_r (794 downto 731) <= data_in(63 downto 0);
                        bits_in_buffer               <= 795;
                    when 732 =>
                        buf_input_r (795 downto 732) <= data_in(63 downto 0);
                        bits_in_buffer               <= 796;
                    when 733 =>
                        buf_input_r (796 downto 733) <= data_in(63 downto 0);
                        bits_in_buffer               <= 797;
                    when 734 =>
                        buf_input_r (797 downto 734) <= data_in(63 downto 0);
                        bits_in_buffer               <= 798;
                    when 735 =>
                        buf_input_r (798 downto 735) <= data_in(63 downto 0);
                        bits_in_buffer               <= 799;
                    when 736 =>
                        buf_input_r (799 downto 736) <= data_in(63 downto 0);
                        bits_in_buffer               <= 800;
                    when 737 =>
                        buf_input_r (800 downto 737) <= data_in(63 downto 0);
                        bits_in_buffer               <= 801;
                    when 738 =>
                        buf_input_r (801 downto 738) <= data_in(63 downto 0);
                        bits_in_buffer               <= 802;
                    when 739 =>
                        buf_input_r (802 downto 739) <= data_in(63 downto 0);
                        bits_in_buffer               <= 803;
                    when 740 =>
                        buf_input_r (803 downto 740) <= data_in(63 downto 0);
                        bits_in_buffer               <= 804;
                    when 741 =>
                        buf_input_r (804 downto 741) <= data_in(63 downto 0);
                        bits_in_buffer               <= 805;
                    when 742 =>
                        buf_input_r (805 downto 742) <= data_in(63 downto 0);
                        bits_in_buffer               <= 806;
                    when 743 =>
                        buf_input_r (806 downto 743) <= data_in(63 downto 0);
                        bits_in_buffer               <= 807;
                    when 744 =>
                        buf_input_r (807 downto 744) <= data_in(63 downto 0);
                        bits_in_buffer               <= 808;
                    when 745 =>
                        buf_input_r (808 downto 745) <= data_in(63 downto 0);
                        bits_in_buffer               <= 809;
                    when 746 =>
                        buf_input_r (809 downto 746) <= data_in(63 downto 0);
                        bits_in_buffer               <= 810;
                    when 747 =>
                        buf_input_r (810 downto 747) <= data_in(63 downto 0);
                        bits_in_buffer               <= 811;
                    when 748 =>
                        buf_input_r (811 downto 748) <= data_in(63 downto 0);
                        bits_in_buffer               <= 812;
                    when 749 =>
                        buf_input_r (812 downto 749) <= data_in(63 downto 0);
                        bits_in_buffer               <= 813;
                    when 750 =>
                        buf_input_r (813 downto 750) <= data_in(63 downto 0);
                        bits_in_buffer               <= 814;
                    when 751 =>
                        buf_input_r (814 downto 751) <= data_in(63 downto 0);
                        bits_in_buffer               <= 815;
                    when 752 =>
                        buf_input_r (815 downto 752) <= data_in(63 downto 0);
                        bits_in_buffer               <= 816;
                    when 753 =>
                        buf_input_r (816 downto 753) <= data_in(63 downto 0);
                        bits_in_buffer               <= 817;
                    when 754 =>
                        buf_input_r (817 downto 754) <= data_in(63 downto 0);
                        bits_in_buffer               <= 818;
                    when 755 =>
                        buf_input_r (818 downto 755) <= data_in(63 downto 0);
                        bits_in_buffer               <= 819;
                    when 756 =>
                        buf_input_r (819 downto 756) <= data_in(63 downto 0);
                        bits_in_buffer               <= 820;
                    when 757 =>
                        buf_input_r (820 downto 757) <= data_in(63 downto 0);
                        bits_in_buffer               <= 821;
                    when 758 =>
                        buf_input_r (821 downto 758) <= data_in(63 downto 0);
                        bits_in_buffer               <= 822;
                    when 759 =>
                        buf_input_r (822 downto 759) <= data_in(63 downto 0);
                        bits_in_buffer               <= 823;
                    when 760 =>
                        buf_input_r (823 downto 760) <= data_in(63 downto 0);
                        bits_in_buffer               <= 824;
                    when 761 =>
                        buf_input_r (824 downto 761) <= data_in(63 downto 0);
                        bits_in_buffer               <= 825;
                    when 762 =>
                        buf_input_r (825 downto 762) <= data_in(63 downto 0);
                        bits_in_buffer               <= 826;
                    when 763 =>
                        buf_input_r (826 downto 763) <= data_in(63 downto 0);
                        bits_in_buffer               <= 827;
                    when 764 =>
                        buf_input_r (827 downto 764) <= data_in(63 downto 0);
                        bits_in_buffer               <= 828;
                    when 765 =>
                        buf_input_r (828 downto 765) <= data_in(63 downto 0);
                        bits_in_buffer               <= 829;
                    when 766 =>
                        buf_input_r (829 downto 766) <= data_in(63 downto 0);
                        bits_in_buffer               <= 830;
                    when 767 =>
                        buf_input_r (830 downto 767) <= data_in(63 downto 0);
                        bits_in_buffer               <= 831;
                    when 768 =>
                        buf_input_r (831 downto 768) <= data_in(63 downto 0);
                        bits_in_buffer               <= 832;
                    when 769 =>
                        buf_input_r (832 downto 769) <= data_in(63 downto 0);
                        bits_in_buffer               <= 833;
                    when 770 =>
                        buf_input_r (833 downto 770) <= data_in(63 downto 0);
                        bits_in_buffer               <= 834;
                    when 771 =>
                        buf_input_r (834 downto 771) <= data_in(63 downto 0);
                        bits_in_buffer               <= 835;
                    when 772 =>
                        buf_input_r (835 downto 772) <= data_in(63 downto 0);
                        bits_in_buffer               <= 836;
                    when 773 =>
                        buf_input_r (836 downto 773) <= data_in(63 downto 0);
                        bits_in_buffer               <= 837;
                    when 774 =>
                        buf_input_r (837 downto 774) <= data_in(63 downto 0);
                        bits_in_buffer               <= 838;
                    when 775 =>
                        buf_input_r (838 downto 775) <= data_in(63 downto 0);
                        bits_in_buffer               <= 839;
                    when 776 =>
                        buf_input_r (839 downto 776) <= data_in(63 downto 0);
                        bits_in_buffer               <= 840;
                    when 777 =>
                        buf_input_r (840 downto 777) <= data_in(63 downto 0);
                        bits_in_buffer               <= 841;
                    when 778 =>
                        buf_input_r (841 downto 778) <= data_in(63 downto 0);
                        bits_in_buffer               <= 842;
                    when 779 =>
                        buf_input_r (842 downto 779) <= data_in(63 downto 0);
                        bits_in_buffer               <= 843;
                    when 780 =>
                        buf_input_r (843 downto 780) <= data_in(63 downto 0);
                        bits_in_buffer               <= 844;
                    when 781 =>
                        buf_input_r (844 downto 781) <= data_in(63 downto 0);
                        bits_in_buffer               <= 845;
                    when 782 =>
                        buf_input_r (845 downto 782) <= data_in(63 downto 0);
                        bits_in_buffer               <= 846;
                    when 783 =>
                        buf_input_r (846 downto 783) <= data_in(63 downto 0);
                        bits_in_buffer               <= 847;
                    when 784 =>
                        buf_input_r (847 downto 784) <= data_in(63 downto 0);
                        bits_in_buffer               <= 848;
                    when 785 =>
                        buf_input_r (848 downto 785) <= data_in(63 downto 0);
                        bits_in_buffer               <= 849;
                    when 786 =>
                        buf_input_r (849 downto 786) <= data_in(63 downto 0);
                        bits_in_buffer               <= 850;
                    when 787 =>
                        buf_input_r (850 downto 787) <= data_in(63 downto 0);
                        bits_in_buffer               <= 851;
                    when 788 =>
                        buf_input_r (851 downto 788) <= data_in(63 downto 0);
                        bits_in_buffer               <= 852;
                    when 789 =>
                        buf_input_r (852 downto 789) <= data_in(63 downto 0);
                        bits_in_buffer               <= 853;
                    when 790 =>
                        buf_input_r (853 downto 790) <= data_in(63 downto 0);
                        bits_in_buffer               <= 854;
                    when 791 =>
                        buf_input_r (854 downto 791) <= data_in(63 downto 0);
                        bits_in_buffer               <= 855;
                    when 792 =>
                        buf_input_r (855 downto 792) <= data_in(63 downto 0);
                        bits_in_buffer               <= 856;
                    when 793 =>
                        buf_input_r (856 downto 793) <= data_in(63 downto 0);
                        bits_in_buffer               <= 857;
                    when 794 =>
                        buf_input_r (857 downto 794) <= data_in(63 downto 0);
                        bits_in_buffer               <= 858;
                    when 795 =>
                        buf_input_r (858 downto 795) <= data_in(63 downto 0);
                        bits_in_buffer               <= 859;
                    when 796 =>
                        buf_input_r (859 downto 796) <= data_in(63 downto 0);
                        bits_in_buffer               <= 860;
                    when 797 =>
                        buf_input_r (860 downto 797) <= data_in(63 downto 0);
                        bits_in_buffer               <= 861;
                    when 798 =>
                        buf_input_r (861 downto 798) <= data_in(63 downto 0);
                        bits_in_buffer               <= 862;
                    when 799 =>
                        buf_input_r (862 downto 799) <= data_in(63 downto 0);
                        bits_in_buffer               <= 863;
                    when 800 =>
                        buf_input_r (863 downto 800) <= data_in(63 downto 0);
                        bits_in_buffer               <= 864;
                    when 801 =>
                        buf_input_r (864 downto 801) <= data_in(63 downto 0);
                        bits_in_buffer               <= 865;
                    when 802 =>
                        buf_input_r (865 downto 802) <= data_in(63 downto 0);
                        bits_in_buffer               <= 866;
                    when 803 =>
                        buf_input_r (866 downto 803) <= data_in(63 downto 0);
                        bits_in_buffer               <= 867;
                    when 804 =>
                        buf_input_r (867 downto 804) <= data_in(63 downto 0);
                        bits_in_buffer               <= 868;
                    when 805 =>
                        buf_input_r (868 downto 805) <= data_in(63 downto 0);
                        bits_in_buffer               <= 869;
                    when 806 =>
                        buf_input_r (869 downto 806) <= data_in(63 downto 0);
                        bits_in_buffer               <= 870;
                    when 807 =>
                        buf_input_r (870 downto 807) <= data_in(63 downto 0);
                        bits_in_buffer               <= 871;
                    when 808 =>
                        buf_input_r (871 downto 808) <= data_in(63 downto 0);
                        bits_in_buffer               <= 872;
                    when 809 =>
                        buf_input_r (872 downto 809) <= data_in(63 downto 0);
                        bits_in_buffer               <= 873;
                    when 810 =>
                        buf_input_r (873 downto 810) <= data_in(63 downto 0);
                        bits_in_buffer               <= 874;
                    when 811 =>
                        buf_input_r (874 downto 811) <= data_in(63 downto 0);
                        bits_in_buffer               <= 875;
                    when 812 =>
                        buf_input_r (875 downto 812) <= data_in(63 downto 0);
                        bits_in_buffer               <= 876;
                    when 813 =>
                        buf_input_r (876 downto 813) <= data_in(63 downto 0);
                        bits_in_buffer               <= 877;
                    when 814 =>
                        buf_input_r (877 downto 814) <= data_in(63 downto 0);
                        bits_in_buffer               <= 878;
                    when 815 =>
                        buf_input_r (878 downto 815) <= data_in(63 downto 0);
                        bits_in_buffer               <= 879;
                    when 816 =>
                        buf_input_r (879 downto 816) <= data_in(63 downto 0);
                        bits_in_buffer               <= 880;
                    when 817 =>
                        buf_input_r (880 downto 817) <= data_in(63 downto 0);
                        bits_in_buffer               <= 881;
                    when 818 =>
                        buf_input_r (881 downto 818) <= data_in(63 downto 0);
                        bits_in_buffer               <= 882;
                    when 819 =>
                        buf_input_r (882 downto 819) <= data_in(63 downto 0);
                        bits_in_buffer               <= 883;
                    when 820 =>
                        buf_input_r (883 downto 820) <= data_in(63 downto 0);
                        bits_in_buffer               <= 884;
                    when 821 =>
                        buf_input_r (884 downto 821) <= data_in(63 downto 0);
                        bits_in_buffer               <= 885;
                    when 822 =>
                        buf_input_r (885 downto 822) <= data_in(63 downto 0);
                        bits_in_buffer               <= 886;
                    when 823 =>
                        buf_input_r (886 downto 823) <= data_in(63 downto 0);
                        bits_in_buffer               <= 887;
                    when 824 =>
                        buf_input_r (887 downto 824) <= data_in(63 downto 0);
                        bits_in_buffer               <= 888;
                    when 825 =>
                        buf_input_r (888 downto 825) <= data_in(63 downto 0);
                        bits_in_buffer               <= 889;
                    when 826 =>
                        buf_input_r (889 downto 826) <= data_in(63 downto 0);
                        bits_in_buffer               <= 890;
                    when 827 =>
                        buf_input_r (890 downto 827) <= data_in(63 downto 0);
                        bits_in_buffer               <= 891;
                    when 828 =>
                        buf_input_r (891 downto 828) <= data_in(63 downto 0);
                        bits_in_buffer               <= 892;
                    when 829 =>
                        buf_input_r (892 downto 829) <= data_in(63 downto 0);
                        bits_in_buffer               <= 893;
                    when 830 =>
                        buf_input_r (893 downto 830) <= data_in(63 downto 0);
                        bits_in_buffer               <= 894;
                    when 831 =>
                        buf_input_r (894 downto 831) <= data_in(63 downto 0);
                        bits_in_buffer               <= 895;
                    when 832 =>
                        buf_input_r (895 downto 832) <= data_in(63 downto 0);
                        bits_in_buffer               <= 896;
                    when 833 =>
                        buf_input_r (896 downto 833) <= data_in(63 downto 0);
                        bits_in_buffer               <= 897;
                    when 834 =>
                        buf_input_r (897 downto 834) <= data_in(63 downto 0);
                        bits_in_buffer               <= 898;
                    when 835 =>
                        buf_input_r (898 downto 835) <= data_in(63 downto 0);
                        bits_in_buffer               <= 899;
                    when 836 =>
                        buf_input_r (899 downto 836) <= data_in(63 downto 0);
                        bits_in_buffer               <= 900;
                    when 837 =>
                        buf_input_r (900 downto 837) <= data_in(63 downto 0);
                        bits_in_buffer               <= 901;
                    when 838 =>
                        buf_input_r (901 downto 838) <= data_in(63 downto 0);
                        bits_in_buffer               <= 902;
                    when 839 =>
                        buf_input_r (902 downto 839) <= data_in(63 downto 0);
                        bits_in_buffer               <= 903;
                    when 840 =>
                        buf_input_r (903 downto 840) <= data_in(63 downto 0);
                        bits_in_buffer               <= 904;
                    when 841 =>
                        buf_input_r (904 downto 841) <= data_in(63 downto 0);
                        bits_in_buffer               <= 905;
                    when 842 =>
                        buf_input_r (905 downto 842) <= data_in(63 downto 0);
                        bits_in_buffer               <= 906;
                    when 843 =>
                        buf_input_r (906 downto 843) <= data_in(63 downto 0);
                        bits_in_buffer               <= 907;
                    when 844 =>
                        buf_input_r (907 downto 844) <= data_in(63 downto 0);
                        bits_in_buffer               <= 908;
                    when 845 =>
                        buf_input_r (908 downto 845) <= data_in(63 downto 0);
                        bits_in_buffer               <= 909;
                    when 846 =>
                        buf_input_r (909 downto 846) <= data_in(63 downto 0);
                        bits_in_buffer               <= 910;
                    when 847 =>
                        buf_input_r (910 downto 847) <= data_in(63 downto 0);
                        bits_in_buffer               <= 911;
                    when 848 =>
                        buf_input_r (911 downto 848) <= data_in(63 downto 0);
                        bits_in_buffer               <= 912;
                    when 849 =>
                        buf_input_r (912 downto 849) <= data_in(63 downto 0);
                        bits_in_buffer               <= 913;
                    when 850 =>
                        buf_input_r (913 downto 850) <= data_in(63 downto 0);
                        bits_in_buffer               <= 914;
                    when 851 =>
                        buf_input_r (914 downto 851) <= data_in(63 downto 0);
                        bits_in_buffer               <= 915;
                    when 852 =>
                        buf_input_r (915 downto 852) <= data_in(63 downto 0);
                        bits_in_buffer               <= 916;
                    when 853 =>
                        buf_input_r (916 downto 853) <= data_in(63 downto 0);
                        bits_in_buffer               <= 917;
                    when 854 =>
                        buf_input_r (917 downto 854) <= data_in(63 downto 0);
                        bits_in_buffer               <= 918;
                    when 855 =>
                        buf_input_r (918 downto 855) <= data_in(63 downto 0);
                        bits_in_buffer               <= 919;
                    when 856 =>
                        buf_input_r (919 downto 856) <= data_in(63 downto 0);
                        bits_in_buffer               <= 920;
                    when 857 =>
                        buf_input_r (920 downto 857) <= data_in(63 downto 0);
                        bits_in_buffer               <= 921;
                    when 858 =>
                        buf_input_r (921 downto 858) <= data_in(63 downto 0);
                        bits_in_buffer               <= 922;
                    when 859 =>
                        buf_input_r (922 downto 859) <= data_in(63 downto 0);
                        bits_in_buffer               <= 923;
                    when 860 =>
                        buf_input_r (923 downto 860) <= data_in(63 downto 0);
                        bits_in_buffer               <= 924;
                    when 861 =>
                        buf_input_r (924 downto 861) <= data_in(63 downto 0);
                        bits_in_buffer               <= 925;
                    when 862 =>
                        buf_input_r (925 downto 862) <= data_in(63 downto 0);
                        bits_in_buffer               <= 926;
                    when 863 =>
                        buf_input_r (926 downto 863) <= data_in(63 downto 0);
                        bits_in_buffer               <= 927;
                    when 864 =>
                        buf_input_r (927 downto 864) <= data_in(63 downto 0);
                        bits_in_buffer               <= 928;
                    when 865 =>
                        buf_input_r (928 downto 865) <= data_in(63 downto 0);
                        bits_in_buffer               <= 929;
                    when 866 =>
                        buf_input_r (929 downto 866) <= data_in(63 downto 0);
                        bits_in_buffer               <= 930;
                    when 867 =>
                        buf_input_r (930 downto 867) <= data_in(63 downto 0);
                        bits_in_buffer               <= 931;
                    when 868 =>
                        buf_input_r (931 downto 868) <= data_in(63 downto 0);
                        bits_in_buffer               <= 932;
                    when 869 =>
                        buf_input_r (932 downto 869) <= data_in(63 downto 0);
                        bits_in_buffer               <= 933;
                    when 870 =>
                        buf_input_r (933 downto 870) <= data_in(63 downto 0);
                        bits_in_buffer               <= 934;
                    when 871 =>
                        buf_input_r (934 downto 871) <= data_in(63 downto 0);
                        bits_in_buffer               <= 935;
                    when 872 =>
                        buf_input_r (935 downto 872) <= data_in(63 downto 0);
                        bits_in_buffer               <= 936;
                    when 873 =>
                        buf_input_r (936 downto 873) <= data_in(63 downto 0);
                        bits_in_buffer               <= 937;
                    when 874 =>
                        buf_input_r (937 downto 874) <= data_in(63 downto 0);
                        bits_in_buffer               <= 938;
                    when 875 =>
                        buf_input_r (938 downto 875) <= data_in(63 downto 0);
                        bits_in_buffer               <= 939;
                    when 876 =>
                        buf_input_r (939 downto 876) <= data_in(63 downto 0);
                        bits_in_buffer               <= 940;
                    when 877 =>
                        buf_input_r (940 downto 877) <= data_in(63 downto 0);
                        bits_in_buffer               <= 941;
                    when 878 =>
                        buf_input_r (941 downto 878) <= data_in(63 downto 0);
                        bits_in_buffer               <= 942;
                    when 879 =>
                        buf_input_r (942 downto 879) <= data_in(63 downto 0);
                        bits_in_buffer               <= 943;
                    when 880 =>
                        buf_input_r (943 downto 880) <= data_in(63 downto 0);
                        bits_in_buffer               <= 944;
                    when 881 =>
                        buf_input_r (944 downto 881) <= data_in(63 downto 0);
                        bits_in_buffer               <= 945;
                    when 882 =>
                        buf_input_r (945 downto 882) <= data_in(63 downto 0);
                        bits_in_buffer               <= 946;
                    when 883 =>
                        buf_input_r (946 downto 883) <= data_in(63 downto 0);
                        bits_in_buffer               <= 947;
                    when 884 =>
                        buf_input_r (947 downto 884) <= data_in(63 downto 0);
                        bits_in_buffer               <= 948;
                    when 885 =>
                        buf_input_r (948 downto 885) <= data_in(63 downto 0);
                        bits_in_buffer               <= 949;
                    when 886 =>
                        buf_input_r (949 downto 886) <= data_in(63 downto 0);
                        bits_in_buffer               <= 950;
                    when 887 =>
                        buf_input_r (950 downto 887) <= data_in(63 downto 0);
                        bits_in_buffer               <= 951;
                    when 888 =>
                        buf_input_r (951 downto 888) <= data_in(63 downto 0);
                        bits_in_buffer               <= 952;
                    when 889 =>
                        buf_input_r (952 downto 889) <= data_in(63 downto 0);
                        bits_in_buffer               <= 953;
                    when 890 =>
                        buf_input_r (953 downto 890) <= data_in(63 downto 0);
                        bits_in_buffer               <= 954;
                    when 891 =>
                        buf_input_r (954 downto 891) <= data_in(63 downto 0);
                        bits_in_buffer               <= 955;
                    when 892 =>
                        buf_input_r (955 downto 892) <= data_in(63 downto 0);
                        bits_in_buffer               <= 956;
                    when 893 =>
                        buf_input_r (956 downto 893) <= data_in(63 downto 0);
                        bits_in_buffer               <= 957;
                    when 894 =>
                        buf_input_r (957 downto 894) <= data_in(63 downto 0);
                        bits_in_buffer               <= 958;
                    when 895 =>
                        buf_input_r (958 downto 895) <= data_in(63 downto 0);
                        bits_in_buffer               <= 959;
                    when 896 =>
                        buf_input_r (959 downto 896) <= data_in(63 downto 0);
                        bits_in_buffer               <= 960;
                    when 897 =>
                        buf_input_r (960 downto 897) <= data_in(63 downto 0);
                        bits_in_buffer               <= 961;
                    when 898 =>
                        buf_input_r (961 downto 898) <= data_in(63 downto 0);
                        bits_in_buffer               <= 962;
                    when 899 =>
                        buf_input_r (962 downto 899) <= data_in(63 downto 0);
                        bits_in_buffer               <= 963;
                    when 900 =>
                        buf_input_r (963 downto 900) <= data_in(63 downto 0);
                        bits_in_buffer               <= 964;
                    when 901 =>
                        buf_input_r (964 downto 901) <= data_in(63 downto 0);
                        bits_in_buffer               <= 965;
                    when 902 =>
                        buf_input_r (965 downto 902) <= data_in(63 downto 0);
                        bits_in_buffer               <= 966;
                    when 903 =>
                        buf_input_r (966 downto 903) <= data_in(63 downto 0);
                        bits_in_buffer               <= 967;
                    when 904 =>
                        buf_input_r (967 downto 904) <= data_in(63 downto 0);
                        bits_in_buffer               <= 968;
                    when 905 =>
                        buf_input_r (968 downto 905) <= data_in(63 downto 0);
                        bits_in_buffer               <= 969;
                    when 906 =>
                        buf_input_r (969 downto 906) <= data_in(63 downto 0);
                        bits_in_buffer               <= 970;
                    when 907 =>
                        buf_input_r (970 downto 907) <= data_in(63 downto 0);
                        bits_in_buffer               <= 971;
                    when 908 =>
                        buf_input_r (971 downto 908) <= data_in(63 downto 0);
                        bits_in_buffer               <= 972;
                    when 909 =>
                        buf_input_r (972 downto 909) <= data_in(63 downto 0);
                        bits_in_buffer               <= 973;
                    when 910 =>
                        buf_input_r (973 downto 910) <= data_in(63 downto 0);
                        bits_in_buffer               <= 974;
                    when 911 =>
                        buf_input_r (974 downto 911) <= data_in(63 downto 0);
                        bits_in_buffer               <= 975;
                    when 912 =>
                        buf_input_r (975 downto 912) <= data_in(63 downto 0);
                        bits_in_buffer               <= 976;
                    when 913 =>
                        buf_input_r (976 downto 913) <= data_in(63 downto 0);
                        bits_in_buffer               <= 977;
                    when 914 =>
                        buf_input_r (977 downto 914) <= data_in(63 downto 0);
                        bits_in_buffer               <= 978;
                    when 915 =>
                        buf_input_r (978 downto 915) <= data_in(63 downto 0);
                        bits_in_buffer               <= 979;
                    when 916 =>
                        buf_input_r (979 downto 916) <= data_in(63 downto 0);
                        bits_in_buffer               <= 980;
                    when 917 =>
                        buf_input_r (980 downto 917) <= data_in(63 downto 0);
                        bits_in_buffer               <= 981;
                    when 918 =>
                        buf_input_r (981 downto 918) <= data_in(63 downto 0);
                        bits_in_buffer               <= 982;
                    when 919 =>
                        buf_input_r (982 downto 919) <= data_in(63 downto 0);
                        bits_in_buffer               <= 983;
                    when 920 =>
                        buf_input_r (983 downto 920) <= data_in(63 downto 0);
                        bits_in_buffer               <= 984;
                    when 921 =>
                        buf_input_r (984 downto 921) <= data_in(63 downto 0);
                        bits_in_buffer               <= 985;
                    when 922 =>
                        buf_input_r (985 downto 922) <= data_in(63 downto 0);
                        bits_in_buffer               <= 986;
                    when 923 =>
                        buf_input_r (986 downto 923) <= data_in(63 downto 0);
                        bits_in_buffer               <= 987;
                    when 924 =>
                        buf_input_r (987 downto 924) <= data_in(63 downto 0);
                        bits_in_buffer               <= 988;
                    when 925 =>
                        buf_input_r (988 downto 925) <= data_in(63 downto 0);
                        bits_in_buffer               <= 989;
                    when 926 =>
                        buf_input_r (989 downto 926) <= data_in(63 downto 0);
                        bits_in_buffer               <= 990;
                    when 927 =>
                        buf_input_r (990 downto 927) <= data_in(63 downto 0);
                        bits_in_buffer               <= 991;
                    when 928 =>
                        buf_input_r (991 downto 928) <= data_in(63 downto 0);
                        bits_in_buffer               <= 992;
                    when 929 =>
                        buf_input_r (992 downto 929) <= data_in(63 downto 0);
                        bits_in_buffer               <= 993;
                    when 930 =>
                        buf_input_r (993 downto 930) <= data_in(63 downto 0);
                        bits_in_buffer               <= 994;
                    when 931 =>
                        buf_input_r (994 downto 931) <= data_in(63 downto 0);
                        bits_in_buffer               <= 995;
                    when 932 =>
                        buf_input_r (995 downto 932) <= data_in(63 downto 0);
                        bits_in_buffer               <= 996;
                    when 933 =>
                        buf_input_r (996 downto 933) <= data_in(63 downto 0);
                        bits_in_buffer               <= 997;
                    when 934 =>
                        buf_input_r (997 downto 934) <= data_in(63 downto 0);
                        bits_in_buffer               <= 998;
                    when 935 =>
                        buf_input_r (998 downto 935) <= data_in(63 downto 0);
                        bits_in_buffer               <= 999;
                    when 936 =>
                        buf_input_r (999 downto 936) <= data_in(63 downto 0);
                        bits_in_buffer               <= 1000;
                    when 937 =>
                        buf_input_r (1000 downto 937) <= data_in(63 downto 0);
                        bits_in_buffer               <= 1001;
                    when 938 =>
                        buf_input_r (1001 downto 938) <= data_in(63 downto 0);
                        bits_in_buffer               <= 1002;
                    when others =>
                end case;
            end if;
        --else
                --out_rdy_r <= '0';
        end if;
    end if;
end process;
end arch_word_expander_64IN_to_1003OUT;