library ieee;
use ieee.std_logic_1164.all;
entity syncalc is
    port(
        in_data     :    in  std_logic_vector(510 downto 0);
        out_data    :    out std_logic_vector(53 downto 0)
);
end entity;

architecture arch of syncalc is
begin
out_data(0)<= in_data(0) xor in_data(9) xor in_data(14) xor in_data(18) xor in_data(19) xor in_data(24) xor in_data(27) xor in_data(28) xor in_data(29) xor in_data(32) xor in_data(34) xor in_data(36) xor in_data(38) xor in_data(39) xor in_data(44) xor in_data(45) xor in_data(47) xor in_data(48) xor in_data(49) xor in_data(50) xor in_data(52) xor in_data(55) xor in_data(56) xor in_data(58) xor in_data(59) xor in_data(60) xor in_data(63) xor in_data(67) xor in_data(69) xor in_data(74) xor in_data(76) xor in_data(78) xor in_data(79) xor in_data(81) xor in_data(84) xor in_data(85) xor in_data(86) xor in_data(87) xor in_data(88) xor in_data(89) xor in_data(91) xor in_data(92) xor in_data(95) xor in_data(98) xor in_data(101) xor in_data(103) xor in_data(104) xor in_data(106) xor in_data(107) xor in_data(108) xor in_data(109) xor in_data(110) xor in_data(111) xor in_data(114) xor in_data(117) xor in_data(118) xor in_data(120) xor in_data(122) xor in_data(125) xor in_data(126) xor in_data(129) xor in_data(130) xor in_data(138) xor in_data(139) xor in_data(143) xor in_data(144) xor in_data(147) xor in_data(149) xor in_data(153) xor in_data(154) xor in_data(156) xor in_data(159) xor in_data(161) xor in_data(162) xor in_data(163) xor in_data(164) xor in_data(165) xor in_data(166) xor in_data(167) xor in_data(169) xor in_data(173) xor in_data(175) xor in_data(176) xor in_data(180) xor in_data(181) xor in_data(182) xor in_data(184) xor in_data(186) xor in_data(187) xor in_data(190) xor in_data(192) xor in_data(193) xor in_data(196) xor in_data(197) xor in_data(198) xor in_data(199) xor in_data(203) xor in_data(204) xor in_data(205) xor in_data(206) xor in_data(207) xor in_data(209) xor in_data(210) xor in_data(211) xor in_data(213) xor in_data(219) xor in_data(220) xor in_data(222) xor in_data(224) xor in_data(225) xor in_data(227) xor in_data(228) xor in_data(230) xor in_data(231) xor in_data(232) xor in_data(234) xor in_data(235) xor in_data(241) xor in_data(243) xor in_data(244) xor in_data(246) xor in_data(248) xor in_data(249) xor in_data(250) xor in_data(251) xor in_data(252) xor in_data(254) xor in_data(256) xor in_data(258) xor in_data(260) xor in_data(267) xor in_data(269) xor in_data(272) xor in_data(274) xor in_data(276) xor in_data(277) xor in_data(278) xor in_data(279) xor in_data(282) xor in_data(284) xor in_data(285) xor in_data(286) xor in_data(288) xor in_data(289) xor in_data(290) xor in_data(297) xor in_data(298) xor in_data(299) xor in_data(302) xor in_data(303) xor in_data(304) xor in_data(306) xor in_data(309) xor in_data(312) xor in_data(313) xor in_data(314) xor in_data(315) xor in_data(317) xor in_data(319) xor in_data(320) xor in_data(321) xor in_data(323) xor in_data(325) xor in_data(329) xor in_data(332) xor in_data(337) xor in_data(338) xor in_data(341) xor in_data(342) xor in_data(343) xor in_data(348) xor in_data(350) xor in_data(351) xor in_data(352) xor in_data(353) xor in_data(355) xor in_data(356) xor in_data(358) xor in_data(359) xor in_data(362) xor in_data(363) xor in_data(365) xor in_data(370) xor in_data(371) xor in_data(372) xor in_data(374) xor in_data(375) xor in_data(376) xor in_data(377) xor in_data(382) xor in_data(383) xor in_data(384) xor in_data(385) xor in_data(386) xor in_data(387) xor in_data(388) xor in_data(389) xor in_data(390) xor in_data(396) xor in_data(397) xor in_data(398) xor in_data(399) xor in_data(401) xor in_data(402) xor in_data(403) xor in_data(404) xor in_data(405) xor in_data(409) xor in_data(411) xor in_data(412) xor in_data(413) xor in_data(416) xor in_data(417) xor in_data(420) xor in_data(426) xor in_data(429) xor in_data(431) xor in_data(434) xor in_data(435) xor in_data(436) xor in_data(438) xor in_data(439) xor in_data(441) xor in_data(445) xor in_data(446) xor in_data(447) xor in_data(448) xor in_data(451) xor in_data(452) xor in_data(453) xor in_data(454) xor in_data(455) xor in_data(458) xor in_data(459) xor in_data(461) xor in_data(462) xor in_data(466) xor in_data(468) xor in_data(470) xor in_data(473) xor in_data(477) xor in_data(478) xor in_data(479) xor in_data(483) xor in_data(484) xor in_data(486) xor in_data(487) xor in_data(489) xor in_data(491) xor in_data(493) xor in_data(494) xor in_data(495) xor in_data(499) xor in_data(502) xor in_data(503) xor in_data(507);

out_data(1)<= in_data(1) xor in_data(10) xor in_data(15) xor in_data(19) xor in_data(20) xor in_data(25) xor in_data(28) xor in_data(29) xor in_data(30) xor in_data(33) xor in_data(35) xor in_data(37) xor in_data(39) xor in_data(40) xor in_data(45) xor in_data(46) xor in_data(48) xor in_data(49) xor in_data(50) xor in_data(51) xor in_data(53) xor in_data(56) xor in_data(57) xor in_data(59) xor in_data(60) xor in_data(61) xor in_data(64) xor in_data(68) xor in_data(70) xor in_data(75) xor in_data(77) xor in_data(79) xor in_data(80) xor in_data(82) xor in_data(85) xor in_data(86) xor in_data(87) xor in_data(88) xor in_data(89) xor in_data(90) xor in_data(92) xor in_data(93) xor in_data(96) xor in_data(99) xor in_data(102) xor in_data(104) xor in_data(105) xor in_data(107) xor in_data(108) xor in_data(109) xor in_data(110) xor in_data(111) xor in_data(112) xor in_data(115) xor in_data(118) xor in_data(119) xor in_data(121) xor in_data(123) xor in_data(126) xor in_data(127) xor in_data(130) xor in_data(131) xor in_data(139) xor in_data(140) xor in_data(144) xor in_data(145) xor in_data(148) xor in_data(150) xor in_data(154) xor in_data(155) xor in_data(157) xor in_data(160) xor in_data(162) xor in_data(163) xor in_data(164) xor in_data(165) xor in_data(166) xor in_data(167) xor in_data(168) xor in_data(170) xor in_data(174) xor in_data(176) xor in_data(177) xor in_data(181) xor in_data(182) xor in_data(183) xor in_data(185) xor in_data(187) xor in_data(188) xor in_data(191) xor in_data(193) xor in_data(194) xor in_data(197) xor in_data(198) xor in_data(199) xor in_data(200) xor in_data(204) xor in_data(205) xor in_data(206) xor in_data(207) xor in_data(208) xor in_data(210) xor in_data(211) xor in_data(212) xor in_data(214) xor in_data(220) xor in_data(221) xor in_data(223) xor in_data(225) xor in_data(226) xor in_data(228) xor in_data(229) xor in_data(231) xor in_data(232) xor in_data(233) xor in_data(235) xor in_data(236) xor in_data(242) xor in_data(244) xor in_data(245) xor in_data(247) xor in_data(249) xor in_data(250) xor in_data(251) xor in_data(252) xor in_data(253) xor in_data(255) xor in_data(257) xor in_data(259) xor in_data(261) xor in_data(268) xor in_data(270) xor in_data(273) xor in_data(275) xor in_data(277) xor in_data(278) xor in_data(279) xor in_data(280) xor in_data(283) xor in_data(285) xor in_data(286) xor in_data(287) xor in_data(289) xor in_data(290) xor in_data(291) xor in_data(298) xor in_data(299) xor in_data(300) xor in_data(303) xor in_data(304) xor in_data(305) xor in_data(307) xor in_data(310) xor in_data(313) xor in_data(314) xor in_data(315) xor in_data(316) xor in_data(318) xor in_data(320) xor in_data(321) xor in_data(322) xor in_data(324) xor in_data(326) xor in_data(330) xor in_data(333) xor in_data(338) xor in_data(339) xor in_data(342) xor in_data(343) xor in_data(344) xor in_data(349) xor in_data(351) xor in_data(352) xor in_data(353) xor in_data(354) xor in_data(356) xor in_data(357) xor in_data(359) xor in_data(360) xor in_data(363) xor in_data(364) xor in_data(366) xor in_data(371) xor in_data(372) xor in_data(373) xor in_data(375) xor in_data(376) xor in_data(377) xor in_data(378) xor in_data(383) xor in_data(384) xor in_data(385) xor in_data(386) xor in_data(387) xor in_data(388) xor in_data(389) xor in_data(390) xor in_data(391) xor in_data(397) xor in_data(398) xor in_data(399) xor in_data(400) xor in_data(402) xor in_data(403) xor in_data(404) xor in_data(405) xor in_data(406) xor in_data(410) xor in_data(412) xor in_data(413) xor in_data(414) xor in_data(417) xor in_data(418) xor in_data(421) xor in_data(427) xor in_data(430) xor in_data(432) xor in_data(435) xor in_data(436) xor in_data(437) xor in_data(439) xor in_data(440) xor in_data(442) xor in_data(446) xor in_data(447) xor in_data(448) xor in_data(449) xor in_data(452) xor in_data(453) xor in_data(454) xor in_data(455) xor in_data(456) xor in_data(459) xor in_data(460) xor in_data(462) xor in_data(463) xor in_data(467) xor in_data(469) xor in_data(471) xor in_data(474) xor in_data(478) xor in_data(479) xor in_data(480) xor in_data(484) xor in_data(485) xor in_data(487) xor in_data(488) xor in_data(490) xor in_data(492) xor in_data(494) xor in_data(495) xor in_data(496) xor in_data(500) xor in_data(503) xor in_data(504) xor in_data(508);

out_data(2)<= in_data(2) xor in_data(11) xor in_data(16) xor in_data(20) xor in_data(21) xor in_data(26) xor in_data(29) xor in_data(30) xor in_data(31) xor in_data(34) xor in_data(36) xor in_data(38) xor in_data(40) xor in_data(41) xor in_data(46) xor in_data(47) xor in_data(49) xor in_data(50) xor in_data(51) xor in_data(52) xor in_data(54) xor in_data(57) xor in_data(58) xor in_data(60) xor in_data(61) xor in_data(62) xor in_data(65) xor in_data(69) xor in_data(71) xor in_data(76) xor in_data(78) xor in_data(80) xor in_data(81) xor in_data(83) xor in_data(86) xor in_data(87) xor in_data(88) xor in_data(89) xor in_data(90) xor in_data(91) xor in_data(93) xor in_data(94) xor in_data(97) xor in_data(100) xor in_data(103) xor in_data(105) xor in_data(106) xor in_data(108) xor in_data(109) xor in_data(110) xor in_data(111) xor in_data(112) xor in_data(113) xor in_data(116) xor in_data(119) xor in_data(120) xor in_data(122) xor in_data(124) xor in_data(127) xor in_data(128) xor in_data(131) xor in_data(132) xor in_data(140) xor in_data(141) xor in_data(145) xor in_data(146) xor in_data(149) xor in_data(151) xor in_data(155) xor in_data(156) xor in_data(158) xor in_data(161) xor in_data(163) xor in_data(164) xor in_data(165) xor in_data(166) xor in_data(167) xor in_data(168) xor in_data(169) xor in_data(171) xor in_data(175) xor in_data(177) xor in_data(178) xor in_data(182) xor in_data(183) xor in_data(184) xor in_data(186) xor in_data(188) xor in_data(189) xor in_data(192) xor in_data(194) xor in_data(195) xor in_data(198) xor in_data(199) xor in_data(200) xor in_data(201) xor in_data(205) xor in_data(206) xor in_data(207) xor in_data(208) xor in_data(209) xor in_data(211) xor in_data(212) xor in_data(213) xor in_data(215) xor in_data(221) xor in_data(222) xor in_data(224) xor in_data(226) xor in_data(227) xor in_data(229) xor in_data(230) xor in_data(232) xor in_data(233) xor in_data(234) xor in_data(236) xor in_data(237) xor in_data(243) xor in_data(245) xor in_data(246) xor in_data(248) xor in_data(250) xor in_data(251) xor in_data(252) xor in_data(253) xor in_data(254) xor in_data(256) xor in_data(258) xor in_data(260) xor in_data(262) xor in_data(269) xor in_data(271) xor in_data(274) xor in_data(276) xor in_data(278) xor in_data(279) xor in_data(280) xor in_data(281) xor in_data(284) xor in_data(286) xor in_data(287) xor in_data(288) xor in_data(290) xor in_data(291) xor in_data(292) xor in_data(299) xor in_data(300) xor in_data(301) xor in_data(304) xor in_data(305) xor in_data(306) xor in_data(308) xor in_data(311) xor in_data(314) xor in_data(315) xor in_data(316) xor in_data(317) xor in_data(319) xor in_data(321) xor in_data(322) xor in_data(323) xor in_data(325) xor in_data(327) xor in_data(331) xor in_data(334) xor in_data(339) xor in_data(340) xor in_data(343) xor in_data(344) xor in_data(345) xor in_data(350) xor in_data(352) xor in_data(353) xor in_data(354) xor in_data(355) xor in_data(357) xor in_data(358) xor in_data(360) xor in_data(361) xor in_data(364) xor in_data(365) xor in_data(367) xor in_data(372) xor in_data(373) xor in_data(374) xor in_data(376) xor in_data(377) xor in_data(378) xor in_data(379) xor in_data(384) xor in_data(385) xor in_data(386) xor in_data(387) xor in_data(388) xor in_data(389) xor in_data(390) xor in_data(391) xor in_data(392) xor in_data(398) xor in_data(399) xor in_data(400) xor in_data(401) xor in_data(403) xor in_data(404) xor in_data(405) xor in_data(406) xor in_data(407) xor in_data(411) xor in_data(413) xor in_data(414) xor in_data(415) xor in_data(418) xor in_data(419) xor in_data(422) xor in_data(428) xor in_data(431) xor in_data(433) xor in_data(436) xor in_data(437) xor in_data(438) xor in_data(440) xor in_data(441) xor in_data(443) xor in_data(447) xor in_data(448) xor in_data(449) xor in_data(450) xor in_data(453) xor in_data(454) xor in_data(455) xor in_data(456) xor in_data(457) xor in_data(460) xor in_data(461) xor in_data(463) xor in_data(464) xor in_data(468) xor in_data(470) xor in_data(472) xor in_data(475) xor in_data(479) xor in_data(480) xor in_data(481) xor in_data(485) xor in_data(486) xor in_data(488) xor in_data(489) xor in_data(491) xor in_data(493) xor in_data(495) xor in_data(496) xor in_data(497) xor in_data(501) xor in_data(504) xor in_data(505) xor in_data(509);

out_data(3)<= in_data(3) xor in_data(12) xor in_data(17) xor in_data(21) xor in_data(22) xor in_data(27) xor in_data(30) xor in_data(31) xor in_data(32) xor in_data(35) xor in_data(37) xor in_data(39) xor in_data(41) xor in_data(42) xor in_data(47) xor in_data(48) xor in_data(50) xor in_data(51) xor in_data(52) xor in_data(53) xor in_data(55) xor in_data(58) xor in_data(59) xor in_data(61) xor in_data(62) xor in_data(63) xor in_data(66) xor in_data(70) xor in_data(72) xor in_data(77) xor in_data(79) xor in_data(81) xor in_data(82) xor in_data(84) xor in_data(87) xor in_data(88) xor in_data(89) xor in_data(90) xor in_data(91) xor in_data(92) xor in_data(94) xor in_data(95) xor in_data(98) xor in_data(101) xor in_data(104) xor in_data(106) xor in_data(107) xor in_data(109) xor in_data(110) xor in_data(111) xor in_data(112) xor in_data(113) xor in_data(114) xor in_data(117) xor in_data(120) xor in_data(121) xor in_data(123) xor in_data(125) xor in_data(128) xor in_data(129) xor in_data(132) xor in_data(133) xor in_data(141) xor in_data(142) xor in_data(146) xor in_data(147) xor in_data(150) xor in_data(152) xor in_data(156) xor in_data(157) xor in_data(159) xor in_data(162) xor in_data(164) xor in_data(165) xor in_data(166) xor in_data(167) xor in_data(168) xor in_data(169) xor in_data(170) xor in_data(172) xor in_data(176) xor in_data(178) xor in_data(179) xor in_data(183) xor in_data(184) xor in_data(185) xor in_data(187) xor in_data(189) xor in_data(190) xor in_data(193) xor in_data(195) xor in_data(196) xor in_data(199) xor in_data(200) xor in_data(201) xor in_data(202) xor in_data(206) xor in_data(207) xor in_data(208) xor in_data(209) xor in_data(210) xor in_data(212) xor in_data(213) xor in_data(214) xor in_data(216) xor in_data(222) xor in_data(223) xor in_data(225) xor in_data(227) xor in_data(228) xor in_data(230) xor in_data(231) xor in_data(233) xor in_data(234) xor in_data(235) xor in_data(237) xor in_data(238) xor in_data(244) xor in_data(246) xor in_data(247) xor in_data(249) xor in_data(251) xor in_data(252) xor in_data(253) xor in_data(254) xor in_data(255) xor in_data(257) xor in_data(259) xor in_data(261) xor in_data(263) xor in_data(270) xor in_data(272) xor in_data(275) xor in_data(277) xor in_data(279) xor in_data(280) xor in_data(281) xor in_data(282) xor in_data(285) xor in_data(287) xor in_data(288) xor in_data(289) xor in_data(291) xor in_data(292) xor in_data(293) xor in_data(300) xor in_data(301) xor in_data(302) xor in_data(305) xor in_data(306) xor in_data(307) xor in_data(309) xor in_data(312) xor in_data(315) xor in_data(316) xor in_data(317) xor in_data(318) xor in_data(320) xor in_data(322) xor in_data(323) xor in_data(324) xor in_data(326) xor in_data(328) xor in_data(332) xor in_data(335) xor in_data(340) xor in_data(341) xor in_data(344) xor in_data(345) xor in_data(346) xor in_data(351) xor in_data(353) xor in_data(354) xor in_data(355) xor in_data(356) xor in_data(358) xor in_data(359) xor in_data(361) xor in_data(362) xor in_data(365) xor in_data(366) xor in_data(368) xor in_data(373) xor in_data(374) xor in_data(375) xor in_data(377) xor in_data(378) xor in_data(379) xor in_data(380) xor in_data(385) xor in_data(386) xor in_data(387) xor in_data(388) xor in_data(389) xor in_data(390) xor in_data(391) xor in_data(392) xor in_data(393) xor in_data(399) xor in_data(400) xor in_data(401) xor in_data(402) xor in_data(404) xor in_data(405) xor in_data(406) xor in_data(407) xor in_data(408) xor in_data(412) xor in_data(414) xor in_data(415) xor in_data(416) xor in_data(419) xor in_data(420) xor in_data(423) xor in_data(429) xor in_data(432) xor in_data(434) xor in_data(437) xor in_data(438) xor in_data(439) xor in_data(441) xor in_data(442) xor in_data(444) xor in_data(448) xor in_data(449) xor in_data(450) xor in_data(451) xor in_data(454) xor in_data(455) xor in_data(456) xor in_data(457) xor in_data(458) xor in_data(461) xor in_data(462) xor in_data(464) xor in_data(465) xor in_data(469) xor in_data(471) xor in_data(473) xor in_data(476) xor in_data(480) xor in_data(481) xor in_data(482) xor in_data(486) xor in_data(487) xor in_data(489) xor in_data(490) xor in_data(492) xor in_data(494) xor in_data(496) xor in_data(497) xor in_data(498) xor in_data(502) xor in_data(505) xor in_data(506) xor in_data(510);

out_data(4)<= in_data(4) xor in_data(9) xor in_data(13) xor in_data(14) xor in_data(19) xor in_data(22) xor in_data(23) xor in_data(24) xor in_data(27) xor in_data(29) xor in_data(31) xor in_data(33) xor in_data(34) xor in_data(39) xor in_data(40) xor in_data(42) xor in_data(43) xor in_data(44) xor in_data(45) xor in_data(47) xor in_data(50) xor in_data(51) xor in_data(53) xor in_data(54) xor in_data(55) xor in_data(58) xor in_data(62) xor in_data(64) xor in_data(69) xor in_data(71) xor in_data(73) xor in_data(74) xor in_data(76) xor in_data(79) xor in_data(80) xor in_data(81) xor in_data(82) xor in_data(83) xor in_data(84) xor in_data(86) xor in_data(87) xor in_data(90) xor in_data(93) xor in_data(96) xor in_data(98) xor in_data(99) xor in_data(101) xor in_data(102) xor in_data(103) xor in_data(104) xor in_data(105) xor in_data(106) xor in_data(109) xor in_data(112) xor in_data(113) xor in_data(115) xor in_data(117) xor in_data(120) xor in_data(121) xor in_data(124) xor in_data(125) xor in_data(133) xor in_data(134) xor in_data(138) xor in_data(139) xor in_data(142) xor in_data(144) xor in_data(148) xor in_data(149) xor in_data(151) xor in_data(154) xor in_data(156) xor in_data(157) xor in_data(158) xor in_data(159) xor in_data(160) xor in_data(161) xor in_data(162) xor in_data(164) xor in_data(168) xor in_data(170) xor in_data(171) xor in_data(175) xor in_data(176) xor in_data(177) xor in_data(179) xor in_data(181) xor in_data(182) xor in_data(185) xor in_data(187) xor in_data(188) xor in_data(191) xor in_data(192) xor in_data(193) xor in_data(194) xor in_data(198) xor in_data(199) xor in_data(200) xor in_data(201) xor in_data(202) xor in_data(204) xor in_data(205) xor in_data(206) xor in_data(208) xor in_data(214) xor in_data(215) xor in_data(217) xor in_data(219) xor in_data(220) xor in_data(222) xor in_data(223) xor in_data(225) xor in_data(226) xor in_data(227) xor in_data(229) xor in_data(230) xor in_data(236) xor in_data(238) xor in_data(239) xor in_data(241) xor in_data(243) xor in_data(244) xor in_data(245) xor in_data(246) xor in_data(247) xor in_data(249) xor in_data(251) xor in_data(253) xor in_data(255) xor in_data(262) xor in_data(264) xor in_data(267) xor in_data(269) xor in_data(271) xor in_data(272) xor in_data(273) xor in_data(274) xor in_data(277) xor in_data(279) xor in_data(280) xor in_data(281) xor in_data(283) xor in_data(284) xor in_data(285) xor in_data(292) xor in_data(293) xor in_data(294) xor in_data(297) xor in_data(298) xor in_data(299) xor in_data(301) xor in_data(304) xor in_data(307) xor in_data(308) xor in_data(309) xor in_data(310) xor in_data(312) xor in_data(314) xor in_data(315) xor in_data(316) xor in_data(318) xor in_data(320) xor in_data(324) xor in_data(327) xor in_data(332) xor in_data(333) xor in_data(336) xor in_data(337) xor in_data(338) xor in_data(343) xor in_data(345) xor in_data(346) xor in_data(347) xor in_data(348) xor in_data(350) xor in_data(351) xor in_data(353) xor in_data(354) xor in_data(357) xor in_data(358) xor in_data(360) xor in_data(365) xor in_data(366) xor in_data(367) xor in_data(369) xor in_data(370) xor in_data(371) xor in_data(372) xor in_data(377) xor in_data(378) xor in_data(379) xor in_data(380) xor in_data(381) xor in_data(382) xor in_data(383) xor in_data(384) xor in_data(385) xor in_data(391) xor in_data(392) xor in_data(393) xor in_data(394) xor in_data(396) xor in_data(397) xor in_data(398) xor in_data(399) xor in_data(400) xor in_data(404) xor in_data(406) xor in_data(407) xor in_data(408) xor in_data(411) xor in_data(412) xor in_data(415) xor in_data(421) xor in_data(424) xor in_data(426) xor in_data(429) xor in_data(430) xor in_data(431) xor in_data(433) xor in_data(434) xor in_data(436) xor in_data(440) xor in_data(441) xor in_data(442) xor in_data(443) xor in_data(446) xor in_data(447) xor in_data(448) xor in_data(449) xor in_data(450) xor in_data(453) xor in_data(454) xor in_data(456) xor in_data(457) xor in_data(461) xor in_data(463) xor in_data(465) xor in_data(468) xor in_data(472) xor in_data(473) xor in_data(474) xor in_data(478) xor in_data(479) xor in_data(481) xor in_data(482) xor in_data(484) xor in_data(486) xor in_data(488) xor in_data(489) xor in_data(490) xor in_data(494) xor in_data(497) xor in_data(498) xor in_data(502) xor in_data(506);

out_data(5)<= in_data(5) xor in_data(10) xor in_data(14) xor in_data(15) xor in_data(20) xor in_data(23) xor in_data(24) xor in_data(25) xor in_data(28) xor in_data(30) xor in_data(32) xor in_data(34) xor in_data(35) xor in_data(40) xor in_data(41) xor in_data(43) xor in_data(44) xor in_data(45) xor in_data(46) xor in_data(48) xor in_data(51) xor in_data(52) xor in_data(54) xor in_data(55) xor in_data(56) xor in_data(59) xor in_data(63) xor in_data(65) xor in_data(70) xor in_data(72) xor in_data(74) xor in_data(75) xor in_data(77) xor in_data(80) xor in_data(81) xor in_data(82) xor in_data(83) xor in_data(84) xor in_data(85) xor in_data(87) xor in_data(88) xor in_data(91) xor in_data(94) xor in_data(97) xor in_data(99) xor in_data(100) xor in_data(102) xor in_data(103) xor in_data(104) xor in_data(105) xor in_data(106) xor in_data(107) xor in_data(110) xor in_data(113) xor in_data(114) xor in_data(116) xor in_data(118) xor in_data(121) xor in_data(122) xor in_data(125) xor in_data(126) xor in_data(134) xor in_data(135) xor in_data(139) xor in_data(140) xor in_data(143) xor in_data(145) xor in_data(149) xor in_data(150) xor in_data(152) xor in_data(155) xor in_data(157) xor in_data(158) xor in_data(159) xor in_data(160) xor in_data(161) xor in_data(162) xor in_data(163) xor in_data(165) xor in_data(169) xor in_data(171) xor in_data(172) xor in_data(176) xor in_data(177) xor in_data(178) xor in_data(180) xor in_data(182) xor in_data(183) xor in_data(186) xor in_data(188) xor in_data(189) xor in_data(192) xor in_data(193) xor in_data(194) xor in_data(195) xor in_data(199) xor in_data(200) xor in_data(201) xor in_data(202) xor in_data(203) xor in_data(205) xor in_data(206) xor in_data(207) xor in_data(209) xor in_data(215) xor in_data(216) xor in_data(218) xor in_data(220) xor in_data(221) xor in_data(223) xor in_data(224) xor in_data(226) xor in_data(227) xor in_data(228) xor in_data(230) xor in_data(231) xor in_data(237) xor in_data(239) xor in_data(240) xor in_data(242) xor in_data(244) xor in_data(245) xor in_data(246) xor in_data(247) xor in_data(248) xor in_data(250) xor in_data(252) xor in_data(254) xor in_data(256) xor in_data(263) xor in_data(265) xor in_data(268) xor in_data(270) xor in_data(272) xor in_data(273) xor in_data(274) xor in_data(275) xor in_data(278) xor in_data(280) xor in_data(281) xor in_data(282) xor in_data(284) xor in_data(285) xor in_data(286) xor in_data(293) xor in_data(294) xor in_data(295) xor in_data(298) xor in_data(299) xor in_data(300) xor in_data(302) xor in_data(305) xor in_data(308) xor in_data(309) xor in_data(310) xor in_data(311) xor in_data(313) xor in_data(315) xor in_data(316) xor in_data(317) xor in_data(319) xor in_data(321) xor in_data(325) xor in_data(328) xor in_data(333) xor in_data(334) xor in_data(337) xor in_data(338) xor in_data(339) xor in_data(344) xor in_data(346) xor in_data(347) xor in_data(348) xor in_data(349) xor in_data(351) xor in_data(352) xor in_data(354) xor in_data(355) xor in_data(358) xor in_data(359) xor in_data(361) xor in_data(366) xor in_data(367) xor in_data(368) xor in_data(370) xor in_data(371) xor in_data(372) xor in_data(373) xor in_data(378) xor in_data(379) xor in_data(380) xor in_data(381) xor in_data(382) xor in_data(383) xor in_data(384) xor in_data(385) xor in_data(386) xor in_data(392) xor in_data(393) xor in_data(394) xor in_data(395) xor in_data(397) xor in_data(398) xor in_data(399) xor in_data(400) xor in_data(401) xor in_data(405) xor in_data(407) xor in_data(408) xor in_data(409) xor in_data(412) xor in_data(413) xor in_data(416) xor in_data(422) xor in_data(425) xor in_data(427) xor in_data(430) xor in_data(431) xor in_data(432) xor in_data(434) xor in_data(435) xor in_data(437) xor in_data(441) xor in_data(442) xor in_data(443) xor in_data(444) xor in_data(447) xor in_data(448) xor in_data(449) xor in_data(450) xor in_data(451) xor in_data(454) xor in_data(455) xor in_data(457) xor in_data(458) xor in_data(462) xor in_data(464) xor in_data(466) xor in_data(469) xor in_data(473) xor in_data(474) xor in_data(475) xor in_data(479) xor in_data(480) xor in_data(482) xor in_data(483) xor in_data(485) xor in_data(487) xor in_data(489) xor in_data(490) xor in_data(491) xor in_data(495) xor in_data(498) xor in_data(499) xor in_data(503) xor in_data(507);

out_data(6)<= in_data(6) xor in_data(11) xor in_data(15) xor in_data(16) xor in_data(21) xor in_data(24) xor in_data(25) xor in_data(26) xor in_data(29) xor in_data(31) xor in_data(33) xor in_data(35) xor in_data(36) xor in_data(41) xor in_data(42) xor in_data(44) xor in_data(45) xor in_data(46) xor in_data(47) xor in_data(49) xor in_data(52) xor in_data(53) xor in_data(55) xor in_data(56) xor in_data(57) xor in_data(60) xor in_data(64) xor in_data(66) xor in_data(71) xor in_data(73) xor in_data(75) xor in_data(76) xor in_data(78) xor in_data(81) xor in_data(82) xor in_data(83) xor in_data(84) xor in_data(85) xor in_data(86) xor in_data(88) xor in_data(89) xor in_data(92) xor in_data(95) xor in_data(98) xor in_data(100) xor in_data(101) xor in_data(103) xor in_data(104) xor in_data(105) xor in_data(106) xor in_data(107) xor in_data(108) xor in_data(111) xor in_data(114) xor in_data(115) xor in_data(117) xor in_data(119) xor in_data(122) xor in_data(123) xor in_data(126) xor in_data(127) xor in_data(135) xor in_data(136) xor in_data(140) xor in_data(141) xor in_data(144) xor in_data(146) xor in_data(150) xor in_data(151) xor in_data(153) xor in_data(156) xor in_data(158) xor in_data(159) xor in_data(160) xor in_data(161) xor in_data(162) xor in_data(163) xor in_data(164) xor in_data(166) xor in_data(170) xor in_data(172) xor in_data(173) xor in_data(177) xor in_data(178) xor in_data(179) xor in_data(181) xor in_data(183) xor in_data(184) xor in_data(187) xor in_data(189) xor in_data(190) xor in_data(193) xor in_data(194) xor in_data(195) xor in_data(196) xor in_data(200) xor in_data(201) xor in_data(202) xor in_data(203) xor in_data(204) xor in_data(206) xor in_data(207) xor in_data(208) xor in_data(210) xor in_data(216) xor in_data(217) xor in_data(219) xor in_data(221) xor in_data(222) xor in_data(224) xor in_data(225) xor in_data(227) xor in_data(228) xor in_data(229) xor in_data(231) xor in_data(232) xor in_data(238) xor in_data(240) xor in_data(241) xor in_data(243) xor in_data(245) xor in_data(246) xor in_data(247) xor in_data(248) xor in_data(249) xor in_data(251) xor in_data(253) xor in_data(255) xor in_data(257) xor in_data(264) xor in_data(266) xor in_data(269) xor in_data(271) xor in_data(273) xor in_data(274) xor in_data(275) xor in_data(276) xor in_data(279) xor in_data(281) xor in_data(282) xor in_data(283) xor in_data(285) xor in_data(286) xor in_data(287) xor in_data(294) xor in_data(295) xor in_data(296) xor in_data(299) xor in_data(300) xor in_data(301) xor in_data(303) xor in_data(306) xor in_data(309) xor in_data(310) xor in_data(311) xor in_data(312) xor in_data(314) xor in_data(316) xor in_data(317) xor in_data(318) xor in_data(320) xor in_data(322) xor in_data(326) xor in_data(329) xor in_data(334) xor in_data(335) xor in_data(338) xor in_data(339) xor in_data(340) xor in_data(345) xor in_data(347) xor in_data(348) xor in_data(349) xor in_data(350) xor in_data(352) xor in_data(353) xor in_data(355) xor in_data(356) xor in_data(359) xor in_data(360) xor in_data(362) xor in_data(367) xor in_data(368) xor in_data(369) xor in_data(371) xor in_data(372) xor in_data(373) xor in_data(374) xor in_data(379) xor in_data(380) xor in_data(381) xor in_data(382) xor in_data(383) xor in_data(384) xor in_data(385) xor in_data(386) xor in_data(387) xor in_data(393) xor in_data(394) xor in_data(395) xor in_data(396) xor in_data(398) xor in_data(399) xor in_data(400) xor in_data(401) xor in_data(402) xor in_data(406) xor in_data(408) xor in_data(409) xor in_data(410) xor in_data(413) xor in_data(414) xor in_data(417) xor in_data(423) xor in_data(426) xor in_data(428) xor in_data(431) xor in_data(432) xor in_data(433) xor in_data(435) xor in_data(436) xor in_data(438) xor in_data(442) xor in_data(443) xor in_data(444) xor in_data(445) xor in_data(448) xor in_data(449) xor in_data(450) xor in_data(451) xor in_data(452) xor in_data(455) xor in_data(456) xor in_data(458) xor in_data(459) xor in_data(463) xor in_data(465) xor in_data(467) xor in_data(470) xor in_data(474) xor in_data(475) xor in_data(476) xor in_data(480) xor in_data(481) xor in_data(483) xor in_data(484) xor in_data(486) xor in_data(488) xor in_data(490) xor in_data(491) xor in_data(492) xor in_data(496) xor in_data(499) xor in_data(500) xor in_data(504) xor in_data(508);

out_data(7)<= in_data(7) xor in_data(12) xor in_data(16) xor in_data(17) xor in_data(22) xor in_data(25) xor in_data(26) xor in_data(27) xor in_data(30) xor in_data(32) xor in_data(34) xor in_data(36) xor in_data(37) xor in_data(42) xor in_data(43) xor in_data(45) xor in_data(46) xor in_data(47) xor in_data(48) xor in_data(50) xor in_data(53) xor in_data(54) xor in_data(56) xor in_data(57) xor in_data(58) xor in_data(61) xor in_data(65) xor in_data(67) xor in_data(72) xor in_data(74) xor in_data(76) xor in_data(77) xor in_data(79) xor in_data(82) xor in_data(83) xor in_data(84) xor in_data(85) xor in_data(86) xor in_data(87) xor in_data(89) xor in_data(90) xor in_data(93) xor in_data(96) xor in_data(99) xor in_data(101) xor in_data(102) xor in_data(104) xor in_data(105) xor in_data(106) xor in_data(107) xor in_data(108) xor in_data(109) xor in_data(112) xor in_data(115) xor in_data(116) xor in_data(118) xor in_data(120) xor in_data(123) xor in_data(124) xor in_data(127) xor in_data(128) xor in_data(136) xor in_data(137) xor in_data(141) xor in_data(142) xor in_data(145) xor in_data(147) xor in_data(151) xor in_data(152) xor in_data(154) xor in_data(157) xor in_data(159) xor in_data(160) xor in_data(161) xor in_data(162) xor in_data(163) xor in_data(164) xor in_data(165) xor in_data(167) xor in_data(171) xor in_data(173) xor in_data(174) xor in_data(178) xor in_data(179) xor in_data(180) xor in_data(182) xor in_data(184) xor in_data(185) xor in_data(188) xor in_data(190) xor in_data(191) xor in_data(194) xor in_data(195) xor in_data(196) xor in_data(197) xor in_data(201) xor in_data(202) xor in_data(203) xor in_data(204) xor in_data(205) xor in_data(207) xor in_data(208) xor in_data(209) xor in_data(211) xor in_data(217) xor in_data(218) xor in_data(220) xor in_data(222) xor in_data(223) xor in_data(225) xor in_data(226) xor in_data(228) xor in_data(229) xor in_data(230) xor in_data(232) xor in_data(233) xor in_data(239) xor in_data(241) xor in_data(242) xor in_data(244) xor in_data(246) xor in_data(247) xor in_data(248) xor in_data(249) xor in_data(250) xor in_data(252) xor in_data(254) xor in_data(256) xor in_data(258) xor in_data(265) xor in_data(267) xor in_data(270) xor in_data(272) xor in_data(274) xor in_data(275) xor in_data(276) xor in_data(277) xor in_data(280) xor in_data(282) xor in_data(283) xor in_data(284) xor in_data(286) xor in_data(287) xor in_data(288) xor in_data(295) xor in_data(296) xor in_data(297) xor in_data(300) xor in_data(301) xor in_data(302) xor in_data(304) xor in_data(307) xor in_data(310) xor in_data(311) xor in_data(312) xor in_data(313) xor in_data(315) xor in_data(317) xor in_data(318) xor in_data(319) xor in_data(321) xor in_data(323) xor in_data(327) xor in_data(330) xor in_data(335) xor in_data(336) xor in_data(339) xor in_data(340) xor in_data(341) xor in_data(346) xor in_data(348) xor in_data(349) xor in_data(350) xor in_data(351) xor in_data(353) xor in_data(354) xor in_data(356) xor in_data(357) xor in_data(360) xor in_data(361) xor in_data(363) xor in_data(368) xor in_data(369) xor in_data(370) xor in_data(372) xor in_data(373) xor in_data(374) xor in_data(375) xor in_data(380) xor in_data(381) xor in_data(382) xor in_data(383) xor in_data(384) xor in_data(385) xor in_data(386) xor in_data(387) xor in_data(388) xor in_data(394) xor in_data(395) xor in_data(396) xor in_data(397) xor in_data(399) xor in_data(400) xor in_data(401) xor in_data(402) xor in_data(403) xor in_data(407) xor in_data(409) xor in_data(410) xor in_data(411) xor in_data(414) xor in_data(415) xor in_data(418) xor in_data(424) xor in_data(427) xor in_data(429) xor in_data(432) xor in_data(433) xor in_data(434) xor in_data(436) xor in_data(437) xor in_data(439) xor in_data(443) xor in_data(444) xor in_data(445) xor in_data(446) xor in_data(449) xor in_data(450) xor in_data(451) xor in_data(452) xor in_data(453) xor in_data(456) xor in_data(457) xor in_data(459) xor in_data(460) xor in_data(464) xor in_data(466) xor in_data(468) xor in_data(471) xor in_data(475) xor in_data(476) xor in_data(477) xor in_data(481) xor in_data(482) xor in_data(484) xor in_data(485) xor in_data(487) xor in_data(489) xor in_data(491) xor in_data(492) xor in_data(493) xor in_data(497) xor in_data(500) xor in_data(501) xor in_data(505) xor in_data(509);

out_data(8)<= in_data(8) xor in_data(13) xor in_data(17) xor in_data(18) xor in_data(23) xor in_data(26) xor in_data(27) xor in_data(28) xor in_data(31) xor in_data(33) xor in_data(35) xor in_data(37) xor in_data(38) xor in_data(43) xor in_data(44) xor in_data(46) xor in_data(47) xor in_data(48) xor in_data(49) xor in_data(51) xor in_data(54) xor in_data(55) xor in_data(57) xor in_data(58) xor in_data(59) xor in_data(62) xor in_data(66) xor in_data(68) xor in_data(73) xor in_data(75) xor in_data(77) xor in_data(78) xor in_data(80) xor in_data(83) xor in_data(84) xor in_data(85) xor in_data(86) xor in_data(87) xor in_data(88) xor in_data(90) xor in_data(91) xor in_data(94) xor in_data(97) xor in_data(100) xor in_data(102) xor in_data(103) xor in_data(105) xor in_data(106) xor in_data(107) xor in_data(108) xor in_data(109) xor in_data(110) xor in_data(113) xor in_data(116) xor in_data(117) xor in_data(119) xor in_data(121) xor in_data(124) xor in_data(125) xor in_data(128) xor in_data(129) xor in_data(137) xor in_data(138) xor in_data(142) xor in_data(143) xor in_data(146) xor in_data(148) xor in_data(152) xor in_data(153) xor in_data(155) xor in_data(158) xor in_data(160) xor in_data(161) xor in_data(162) xor in_data(163) xor in_data(164) xor in_data(165) xor in_data(166) xor in_data(168) xor in_data(172) xor in_data(174) xor in_data(175) xor in_data(179) xor in_data(180) xor in_data(181) xor in_data(183) xor in_data(185) xor in_data(186) xor in_data(189) xor in_data(191) xor in_data(192) xor in_data(195) xor in_data(196) xor in_data(197) xor in_data(198) xor in_data(202) xor in_data(203) xor in_data(204) xor in_data(205) xor in_data(206) xor in_data(208) xor in_data(209) xor in_data(210) xor in_data(212) xor in_data(218) xor in_data(219) xor in_data(221) xor in_data(223) xor in_data(224) xor in_data(226) xor in_data(227) xor in_data(229) xor in_data(230) xor in_data(231) xor in_data(233) xor in_data(234) xor in_data(240) xor in_data(242) xor in_data(243) xor in_data(245) xor in_data(247) xor in_data(248) xor in_data(249) xor in_data(250) xor in_data(251) xor in_data(253) xor in_data(255) xor in_data(257) xor in_data(259) xor in_data(266) xor in_data(268) xor in_data(271) xor in_data(273) xor in_data(275) xor in_data(276) xor in_data(277) xor in_data(278) xor in_data(281) xor in_data(283) xor in_data(284) xor in_data(285) xor in_data(287) xor in_data(288) xor in_data(289) xor in_data(296) xor in_data(297) xor in_data(298) xor in_data(301) xor in_data(302) xor in_data(303) xor in_data(305) xor in_data(308) xor in_data(311) xor in_data(312) xor in_data(313) xor in_data(314) xor in_data(316) xor in_data(318) xor in_data(319) xor in_data(320) xor in_data(322) xor in_data(324) xor in_data(328) xor in_data(331) xor in_data(336) xor in_data(337) xor in_data(340) xor in_data(341) xor in_data(342) xor in_data(347) xor in_data(349) xor in_data(350) xor in_data(351) xor in_data(352) xor in_data(354) xor in_data(355) xor in_data(357) xor in_data(358) xor in_data(361) xor in_data(362) xor in_data(364) xor in_data(369) xor in_data(370) xor in_data(371) xor in_data(373) xor in_data(374) xor in_data(375) xor in_data(376) xor in_data(381) xor in_data(382) xor in_data(383) xor in_data(384) xor in_data(385) xor in_data(386) xor in_data(387) xor in_data(388) xor in_data(389) xor in_data(395) xor in_data(396) xor in_data(397) xor in_data(398) xor in_data(400) xor in_data(401) xor in_data(402) xor in_data(403) xor in_data(404) xor in_data(408) xor in_data(410) xor in_data(411) xor in_data(412) xor in_data(415) xor in_data(416) xor in_data(419) xor in_data(425) xor in_data(428) xor in_data(430) xor in_data(433) xor in_data(434) xor in_data(435) xor in_data(437) xor in_data(438) xor in_data(440) xor in_data(444) xor in_data(445) xor in_data(446) xor in_data(447) xor in_data(450) xor in_data(451) xor in_data(452) xor in_data(453) xor in_data(454) xor in_data(457) xor in_data(458) xor in_data(460) xor in_data(461) xor in_data(465) xor in_data(467) xor in_data(469) xor in_data(472) xor in_data(476) xor in_data(477) xor in_data(478) xor in_data(482) xor in_data(483) xor in_data(485) xor in_data(486) xor in_data(488) xor in_data(490) xor in_data(492) xor in_data(493) xor in_data(494) xor in_data(498) xor in_data(501) xor in_data(502) xor in_data(506) xor in_data(510);

out_data(9)<='0';

out_data(10)<='0';

out_data(11)<='0';

out_data(12)<='0';

out_data(13)<='0';

out_data(14)<='0';

out_data(15)<='0';

out_data(16)<='0';

out_data(17)<='0';

out_data(18)<= in_data(0) xor in_data(3) xor in_data(6) xor in_data(8) xor in_data(9) xor in_data(12) xor in_data(13) xor in_data(15) xor in_data(16) xor in_data(20) xor in_data(21) xor in_data(23) xor in_data(26) xor in_data(27) xor in_data(28) xor in_data(29) xor in_data(36) xor in_data(37) xor in_data(38) xor in_data(39) xor in_data(40) xor in_data(42) xor in_data(43) xor in_data(46) xor in_data(48) xor in_data(49) xor in_data(51) xor in_data(52) xor in_data(53) xor in_data(54) xor in_data(55) xor in_data(60) xor in_data(62) xor in_data(64) xor in_data(66) xor in_data(68) xor in_data(69) xor in_data(70) xor in_data(71) xor in_data(73) xor in_data(74) xor in_data(75) xor in_data(76) xor in_data(77) xor in_data(78) xor in_data(81) xor in_data(82) xor in_data(83) xor in_data(84) xor in_data(86) xor in_data(89) xor in_data(92) xor in_data(93) xor in_data(94) xor in_data(95) xor in_data(96) xor in_data(99) xor in_data(101) xor in_data(102) xor in_data(103) xor in_data(104) xor in_data(105) xor in_data(107) xor in_data(114) xor in_data(116) xor in_data(117) xor in_data(121) xor in_data(124) xor in_data(125) xor in_data(128) xor in_data(129) xor in_data(130) xor in_data(132) xor in_data(133) xor in_data(134) xor in_data(135) xor in_data(137) xor in_data(139) xor in_data(140) xor in_data(142) xor in_data(143) xor in_data(145) xor in_data(146) xor in_data(147) xor in_data(149) xor in_data(151) xor in_data(153) xor in_data(154) xor in_data(156) xor in_data(159) xor in_data(161) xor in_data(162) xor in_data(163) xor in_data(165) xor in_data(169) xor in_data(175) xor in_data(180) xor in_data(181) xor in_data(183) xor in_data(185) xor in_data(186) xor in_data(187) xor in_data(189) xor in_data(190) xor in_data(195) xor in_data(199) xor in_data(200) xor in_data(201) xor in_data(202) xor in_data(203) xor in_data(204) xor in_data(205) xor in_data(206) xor in_data(207) xor in_data(211) xor in_data(212) xor in_data(218) xor in_data(220) xor in_data(224) xor in_data(225) xor in_data(226) xor in_data(228) xor in_data(229) xor in_data(231) xor in_data(236) xor in_data(238) xor in_data(239) xor in_data(240) xor in_data(245) xor in_data(246) xor in_data(247) xor in_data(253) xor in_data(254) xor in_data(255) xor in_data(257) xor in_data(260) xor in_data(261) xor in_data(263) xor in_data(265) xor in_data(267) xor in_data(270) xor in_data(271) xor in_data(275) xor in_data(276) xor in_data(277) xor in_data(278) xor in_data(280) xor in_data(281) xor in_data(283) xor in_data(284) xor in_data(287) xor in_data(288) xor in_data(289) xor in_data(290) xor in_data(291) xor in_data(292) xor in_data(294) xor in_data(295) xor in_data(296) xor in_data(298) xor in_data(299) xor in_data(300) xor in_data(303) xor in_data(304) xor in_data(305) xor in_data(308) xor in_data(309) xor in_data(314) xor in_data(315) xor in_data(319) xor in_data(321) xor in_data(322) xor in_data(323) xor in_data(324) xor in_data(327) xor in_data(328) xor in_data(330) xor in_data(334) xor in_data(335) xor in_data(338) xor in_data(347) xor in_data(350) xor in_data(352) xor in_data(357) xor in_data(358) xor in_data(359) xor in_data(360) xor in_data(363) xor in_data(366) xor in_data(367) xor in_data(369) xor in_data(370) xor in_data(371) xor in_data(375) xor in_data(376) xor in_data(377) xor in_data(380) xor in_data(384) xor in_data(387) xor in_data(392) xor in_data(395) xor in_data(396) xor in_data(397) xor in_data(399) xor in_data(401) xor in_data(402) xor in_data(403) xor in_data(404) xor in_data(405) xor in_data(406) xor in_data(407) xor in_data(409) xor in_data(411) xor in_data(414) xor in_data(418) xor in_data(419) xor in_data(421) xor in_data(422) xor in_data(424) xor in_data(426) xor in_data(432) xor in_data(433) xor in_data(436) xor in_data(437) xor in_data(440) xor in_data(442) xor in_data(445) xor in_data(447) xor in_data(449) xor in_data(453) xor in_data(455) xor in_data(458) xor in_data(459) xor in_data(460) xor in_data(464) xor in_data(466) xor in_data(468) xor in_data(469) xor in_data(470) xor in_data(473) xor in_data(475) xor in_data(477) xor in_data(478) xor in_data(486) xor in_data(487) xor in_data(489) xor in_data(490) xor in_data(491) xor in_data(492) xor in_data(496) xor in_data(500) xor in_data(502) xor in_data(503) xor in_data(505) xor in_data(507) xor in_data(508);

out_data(19)<= in_data(5) xor in_data(10) xor in_data(11) xor in_data(13) xor in_data(15) xor in_data(16) xor in_data(17) xor in_data(19) xor in_data(20) xor in_data(25) xor in_data(29) xor in_data(30) xor in_data(31) xor in_data(32) xor in_data(33) xor in_data(34) xor in_data(35) xor in_data(36) xor in_data(37) xor in_data(41) xor in_data(42) xor in_data(48) xor in_data(50) xor in_data(54) xor in_data(55) xor in_data(56) xor in_data(58) xor in_data(59) xor in_data(61) xor in_data(66) xor in_data(68) xor in_data(69) xor in_data(70) xor in_data(75) xor in_data(76) xor in_data(77) xor in_data(83) xor in_data(84) xor in_data(85) xor in_data(87) xor in_data(90) xor in_data(91) xor in_data(93) xor in_data(95) xor in_data(97) xor in_data(100) xor in_data(101) xor in_data(105) xor in_data(106) xor in_data(107) xor in_data(108) xor in_data(110) xor in_data(111) xor in_data(113) xor in_data(114) xor in_data(117) xor in_data(118) xor in_data(119) xor in_data(120) xor in_data(121) xor in_data(122) xor in_data(124) xor in_data(125) xor in_data(126) xor in_data(128) xor in_data(129) xor in_data(130) xor in_data(133) xor in_data(134) xor in_data(135) xor in_data(138) xor in_data(139) xor in_data(144) xor in_data(145) xor in_data(149) xor in_data(151) xor in_data(152) xor in_data(153) xor in_data(154) xor in_data(157) xor in_data(158) xor in_data(160) xor in_data(164) xor in_data(165) xor in_data(168) xor in_data(177) xor in_data(180) xor in_data(182) xor in_data(187) xor in_data(188) xor in_data(189) xor in_data(190) xor in_data(193) xor in_data(196) xor in_data(197) xor in_data(199) xor in_data(200) xor in_data(201) xor in_data(205) xor in_data(206) xor in_data(207) xor in_data(210) xor in_data(214) xor in_data(217) xor in_data(222) xor in_data(225) xor in_data(226) xor in_data(227) xor in_data(229) xor in_data(231) xor in_data(232) xor in_data(233) xor in_data(234) xor in_data(235) xor in_data(236) xor in_data(237) xor in_data(239) xor in_data(241) xor in_data(244) xor in_data(248) xor in_data(249) xor in_data(251) xor in_data(252) xor in_data(254) xor in_data(256) xor in_data(262) xor in_data(263) xor in_data(266) xor in_data(267) xor in_data(270) xor in_data(272) xor in_data(275) xor in_data(277) xor in_data(279) xor in_data(283) xor in_data(285) xor in_data(288) xor in_data(289) xor in_data(290) xor in_data(294) xor in_data(296) xor in_data(298) xor in_data(299) xor in_data(300) xor in_data(303) xor in_data(305) xor in_data(307) xor in_data(308) xor in_data(316) xor in_data(317) xor in_data(319) xor in_data(320) xor in_data(321) xor in_data(322) xor in_data(326) xor in_data(330) xor in_data(332) xor in_data(333) xor in_data(335) xor in_data(337) xor in_data(338) xor in_data(341) xor in_data(344) xor in_data(347) xor in_data(349) xor in_data(350) xor in_data(353) xor in_data(354) xor in_data(356) xor in_data(357) xor in_data(361) xor in_data(362) xor in_data(364) xor in_data(367) xor in_data(368) xor in_data(369) xor in_data(370) xor in_data(377) xor in_data(378) xor in_data(379) xor in_data(380) xor in_data(381) xor in_data(383) xor in_data(384) xor in_data(387) xor in_data(389) xor in_data(390) xor in_data(392) xor in_data(393) xor in_data(394) xor in_data(395) xor in_data(396) xor in_data(401) xor in_data(403) xor in_data(405) xor in_data(407) xor in_data(409) xor in_data(410) xor in_data(411) xor in_data(412) xor in_data(414) xor in_data(415) xor in_data(416) xor in_data(417) xor in_data(418) xor in_data(419) xor in_data(422) xor in_data(423) xor in_data(424) xor in_data(425) xor in_data(427) xor in_data(430) xor in_data(433) xor in_data(434) xor in_data(435) xor in_data(436) xor in_data(437) xor in_data(440) xor in_data(442) xor in_data(443) xor in_data(444) xor in_data(445) xor in_data(446) xor in_data(448) xor in_data(455) xor in_data(457) xor in_data(458) xor in_data(462) xor in_data(465) xor in_data(466) xor in_data(469) xor in_data(470) xor in_data(471) xor in_data(473) xor in_data(474) xor in_data(475) xor in_data(476) xor in_data(478) xor in_data(480) xor in_data(481) xor in_data(483) xor in_data(484) xor in_data(486) xor in_data(487) xor in_data(488) xor in_data(490) xor in_data(492) xor in_data(494) xor in_data(495) xor in_data(497) xor in_data(500) xor in_data(502) xor in_data(503) xor in_data(504) xor in_data(506) xor in_data(510);

out_data(20)<= in_data(7) xor in_data(10) xor in_data(12) xor in_data(17) xor in_data(18) xor in_data(19) xor in_data(20) xor in_data(23) xor in_data(26) xor in_data(27) xor in_data(29) xor in_data(30) xor in_data(31) xor in_data(35) xor in_data(36) xor in_data(37) xor in_data(40) xor in_data(44) xor in_data(47) xor in_data(52) xor in_data(55) xor in_data(56) xor in_data(57) xor in_data(59) xor in_data(61) xor in_data(62) xor in_data(63) xor in_data(64) xor in_data(65) xor in_data(66) xor in_data(67) xor in_data(69) xor in_data(71) xor in_data(74) xor in_data(78) xor in_data(79) xor in_data(81) xor in_data(82) xor in_data(84) xor in_data(86) xor in_data(92) xor in_data(93) xor in_data(96) xor in_data(97) xor in_data(100) xor in_data(102) xor in_data(105) xor in_data(107) xor in_data(109) xor in_data(113) xor in_data(115) xor in_data(118) xor in_data(119) xor in_data(120) xor in_data(124) xor in_data(126) xor in_data(128) xor in_data(129) xor in_data(130) xor in_data(133) xor in_data(135) xor in_data(137) xor in_data(138) xor in_data(146) xor in_data(147) xor in_data(149) xor in_data(150) xor in_data(151) xor in_data(152) xor in_data(156) xor in_data(160) xor in_data(162) xor in_data(163) xor in_data(165) xor in_data(167) xor in_data(168) xor in_data(171) xor in_data(174) xor in_data(177) xor in_data(179) xor in_data(180) xor in_data(183) xor in_data(184) xor in_data(186) xor in_data(187) xor in_data(191) xor in_data(192) xor in_data(194) xor in_data(197) xor in_data(198) xor in_data(199) xor in_data(200) xor in_data(207) xor in_data(208) xor in_data(209) xor in_data(210) xor in_data(211) xor in_data(213) xor in_data(214) xor in_data(217) xor in_data(219) xor in_data(220) xor in_data(222) xor in_data(223) xor in_data(224) xor in_data(225) xor in_data(226) xor in_data(231) xor in_data(233) xor in_data(235) xor in_data(237) xor in_data(239) xor in_data(240) xor in_data(241) xor in_data(242) xor in_data(244) xor in_data(245) xor in_data(246) xor in_data(247) xor in_data(248) xor in_data(249) xor in_data(252) xor in_data(253) xor in_data(254) xor in_data(255) xor in_data(257) xor in_data(260) xor in_data(263) xor in_data(264) xor in_data(265) xor in_data(266) xor in_data(267) xor in_data(270) xor in_data(272) xor in_data(273) xor in_data(274) xor in_data(275) xor in_data(276) xor in_data(278) xor in_data(285) xor in_data(287) xor in_data(288) xor in_data(292) xor in_data(295) xor in_data(296) xor in_data(299) xor in_data(300) xor in_data(301) xor in_data(303) xor in_data(304) xor in_data(305) xor in_data(306) xor in_data(308) xor in_data(310) xor in_data(311) xor in_data(313) xor in_data(314) xor in_data(316) xor in_data(317) xor in_data(318) xor in_data(320) xor in_data(322) xor in_data(324) xor in_data(325) xor in_data(327) xor in_data(330) xor in_data(332) xor in_data(333) xor in_data(334) xor in_data(336) xor in_data(340) xor in_data(346) xor in_data(351) xor in_data(352) xor in_data(354) xor in_data(356) xor in_data(357) xor in_data(358) xor in_data(360) xor in_data(361) xor in_data(366) xor in_data(370) xor in_data(371) xor in_data(372) xor in_data(373) xor in_data(374) xor in_data(375) xor in_data(376) xor in_data(377) xor in_data(378) xor in_data(382) xor in_data(383) xor in_data(389) xor in_data(391) xor in_data(395) xor in_data(396) xor in_data(397) xor in_data(399) xor in_data(400) xor in_data(402) xor in_data(407) xor in_data(409) xor in_data(410) xor in_data(411) xor in_data(416) xor in_data(417) xor in_data(418) xor in_data(424) xor in_data(425) xor in_data(426) xor in_data(428) xor in_data(431) xor in_data(432) xor in_data(434) xor in_data(436) xor in_data(438) xor in_data(441) xor in_data(442) xor in_data(446) xor in_data(447) xor in_data(448) xor in_data(449) xor in_data(451) xor in_data(452) xor in_data(454) xor in_data(455) xor in_data(458) xor in_data(459) xor in_data(460) xor in_data(461) xor in_data(462) xor in_data(463) xor in_data(465) xor in_data(466) xor in_data(467) xor in_data(469) xor in_data(470) xor in_data(471) xor in_data(474) xor in_data(475) xor in_data(476) xor in_data(479) xor in_data(480) xor in_data(485) xor in_data(486) xor in_data(490) xor in_data(492) xor in_data(493) xor in_data(494) xor in_data(495) xor in_data(498) xor in_data(499) xor in_data(501) xor in_data(505) xor in_data(506) xor in_data(509);

out_data(21)<= in_data(1) xor in_data(4) xor in_data(7) xor in_data(9) xor in_data(10) xor in_data(13) xor in_data(14) xor in_data(16) xor in_data(17) xor in_data(21) xor in_data(22) xor in_data(24) xor in_data(27) xor in_data(28) xor in_data(29) xor in_data(30) xor in_data(37) xor in_data(38) xor in_data(39) xor in_data(40) xor in_data(41) xor in_data(43) xor in_data(44) xor in_data(47) xor in_data(49) xor in_data(50) xor in_data(52) xor in_data(53) xor in_data(54) xor in_data(55) xor in_data(56) xor in_data(61) xor in_data(63) xor in_data(65) xor in_data(67) xor in_data(69) xor in_data(70) xor in_data(71) xor in_data(72) xor in_data(74) xor in_data(75) xor in_data(76) xor in_data(77) xor in_data(78) xor in_data(79) xor in_data(82) xor in_data(83) xor in_data(84) xor in_data(85) xor in_data(87) xor in_data(90) xor in_data(93) xor in_data(94) xor in_data(95) xor in_data(96) xor in_data(97) xor in_data(100) xor in_data(102) xor in_data(103) xor in_data(104) xor in_data(105) xor in_data(106) xor in_data(108) xor in_data(115) xor in_data(117) xor in_data(118) xor in_data(122) xor in_data(125) xor in_data(126) xor in_data(129) xor in_data(130) xor in_data(131) xor in_data(133) xor in_data(134) xor in_data(135) xor in_data(136) xor in_data(138) xor in_data(140) xor in_data(141) xor in_data(143) xor in_data(144) xor in_data(146) xor in_data(147) xor in_data(148) xor in_data(150) xor in_data(152) xor in_data(154) xor in_data(155) xor in_data(157) xor in_data(160) xor in_data(162) xor in_data(163) xor in_data(164) xor in_data(166) xor in_data(170) xor in_data(176) xor in_data(181) xor in_data(182) xor in_data(184) xor in_data(186) xor in_data(187) xor in_data(188) xor in_data(190) xor in_data(191) xor in_data(196) xor in_data(200) xor in_data(201) xor in_data(202) xor in_data(203) xor in_data(204) xor in_data(205) xor in_data(206) xor in_data(207) xor in_data(208) xor in_data(212) xor in_data(213) xor in_data(219) xor in_data(221) xor in_data(225) xor in_data(226) xor in_data(227) xor in_data(229) xor in_data(230) xor in_data(232) xor in_data(237) xor in_data(239) xor in_data(240) xor in_data(241) xor in_data(246) xor in_data(247) xor in_data(248) xor in_data(254) xor in_data(255) xor in_data(256) xor in_data(258) xor in_data(261) xor in_data(262) xor in_data(264) xor in_data(266) xor in_data(268) xor in_data(271) xor in_data(272) xor in_data(276) xor in_data(277) xor in_data(278) xor in_data(279) xor in_data(281) xor in_data(282) xor in_data(284) xor in_data(285) xor in_data(288) xor in_data(289) xor in_data(290) xor in_data(291) xor in_data(292) xor in_data(293) xor in_data(295) xor in_data(296) xor in_data(297) xor in_data(299) xor in_data(300) xor in_data(301) xor in_data(304) xor in_data(305) xor in_data(306) xor in_data(309) xor in_data(310) xor in_data(315) xor in_data(316) xor in_data(320) xor in_data(322) xor in_data(323) xor in_data(324) xor in_data(325) xor in_data(328) xor in_data(329) xor in_data(331) xor in_data(335) xor in_data(336) xor in_data(339) xor in_data(348) xor in_data(351) xor in_data(353) xor in_data(358) xor in_data(359) xor in_data(360) xor in_data(361) xor in_data(364) xor in_data(367) xor in_data(368) xor in_data(370) xor in_data(371) xor in_data(372) xor in_data(376) xor in_data(377) xor in_data(378) xor in_data(381) xor in_data(385) xor in_data(388) xor in_data(393) xor in_data(396) xor in_data(397) xor in_data(398) xor in_data(400) xor in_data(402) xor in_data(403) xor in_data(404) xor in_data(405) xor in_data(406) xor in_data(407) xor in_data(408) xor in_data(410) xor in_data(412) xor in_data(415) xor in_data(419) xor in_data(420) xor in_data(422) xor in_data(423) xor in_data(425) xor in_data(427) xor in_data(433) xor in_data(434) xor in_data(437) xor in_data(438) xor in_data(441) xor in_data(443) xor in_data(446) xor in_data(448) xor in_data(450) xor in_data(454) xor in_data(456) xor in_data(459) xor in_data(460) xor in_data(461) xor in_data(465) xor in_data(467) xor in_data(469) xor in_data(470) xor in_data(471) xor in_data(474) xor in_data(476) xor in_data(478) xor in_data(479) xor in_data(487) xor in_data(488) xor in_data(490) xor in_data(491) xor in_data(492) xor in_data(493) xor in_data(497) xor in_data(501) xor in_data(503) xor in_data(504) xor in_data(506) xor in_data(508) xor in_data(509);

out_data(22)<= in_data(3) xor in_data(8) xor in_data(9) xor in_data(11) xor in_data(13) xor in_data(14) xor in_data(15) xor in_data(17) xor in_data(18) xor in_data(23) xor in_data(27) xor in_data(28) xor in_data(29) xor in_data(30) xor in_data(31) xor in_data(32) xor in_data(33) xor in_data(34) xor in_data(35) xor in_data(39) xor in_data(40) xor in_data(46) xor in_data(48) xor in_data(52) xor in_data(53) xor in_data(54) xor in_data(56) xor in_data(57) xor in_data(59) xor in_data(64) xor in_data(66) xor in_data(67) xor in_data(68) xor in_data(73) xor in_data(74) xor in_data(75) xor in_data(81) xor in_data(82) xor in_data(83) xor in_data(85) xor in_data(88) xor in_data(89) xor in_data(91) xor in_data(93) xor in_data(95) xor in_data(98) xor in_data(99) xor in_data(103) xor in_data(104) xor in_data(105) xor in_data(106) xor in_data(108) xor in_data(109) xor in_data(111) xor in_data(112) xor in_data(115) xor in_data(116) xor in_data(117) xor in_data(118) xor in_data(119) xor in_data(120) xor in_data(122) xor in_data(123) xor in_data(124) xor in_data(126) xor in_data(127) xor in_data(128) xor in_data(131) xor in_data(132) xor in_data(133) xor in_data(136) xor in_data(137) xor in_data(142) xor in_data(143) xor in_data(147) xor in_data(149) xor in_data(150) xor in_data(151) xor in_data(152) xor in_data(155) xor in_data(156) xor in_data(158) xor in_data(162) xor in_data(163) xor in_data(166) xor in_data(175) xor in_data(178) xor in_data(180) xor in_data(185) xor in_data(186) xor in_data(187) xor in_data(188) xor in_data(191) xor in_data(194) xor in_data(195) xor in_data(197) xor in_data(198) xor in_data(199) xor in_data(203) xor in_data(204) xor in_data(205) xor in_data(208) xor in_data(212) xor in_data(215) xor in_data(220) xor in_data(223) xor in_data(224) xor in_data(225) xor in_data(227) xor in_data(229) xor in_data(230) xor in_data(231) xor in_data(232) xor in_data(233) xor in_data(234) xor in_data(235) xor in_data(237) xor in_data(239) xor in_data(242) xor in_data(246) xor in_data(247) xor in_data(249) xor in_data(250) xor in_data(252) xor in_data(254) xor in_data(260) xor in_data(261) xor in_data(264) xor in_data(265) xor in_data(268) xor in_data(270) xor in_data(273) xor in_data(275) xor in_data(277) xor in_data(281) xor in_data(283) xor in_data(286) xor in_data(287) xor in_data(288) xor in_data(292) xor in_data(294) xor in_data(296) xor in_data(297) xor in_data(298) xor in_data(301) xor in_data(303) xor in_data(305) xor in_data(306) xor in_data(314) xor in_data(315) xor in_data(317) xor in_data(318) xor in_data(319) xor in_data(320) xor in_data(324) xor in_data(328) xor in_data(330) xor in_data(331) xor in_data(333) xor in_data(335) xor in_data(336) xor in_data(339) xor in_data(342) xor in_data(345) xor in_data(347) xor in_data(348) xor in_data(351) xor in_data(352) xor in_data(354) xor in_data(355) xor in_data(359) xor in_data(360) xor in_data(362) xor in_data(365) xor in_data(366) xor in_data(367) xor in_data(368) xor in_data(375) xor in_data(376) xor in_data(377) xor in_data(378) xor in_data(379) xor in_data(381) xor in_data(382) xor in_data(385) xor in_data(387) xor in_data(388) xor in_data(390) xor in_data(391) xor in_data(392) xor in_data(393) xor in_data(394) xor in_data(399) xor in_data(401) xor in_data(403) xor in_data(405) xor in_data(407) xor in_data(408) xor in_data(409) xor in_data(410) xor in_data(412) xor in_data(413) xor in_data(414) xor in_data(415) xor in_data(416) xor in_data(417) xor in_data(420) xor in_data(421) xor in_data(422) xor in_data(423) xor in_data(425) xor in_data(428) xor in_data(431) xor in_data(432) xor in_data(433) xor in_data(434) xor in_data(435) xor in_data(438) xor in_data(440) xor in_data(441) xor in_data(442) xor in_data(443) xor in_data(444) xor in_data(446) xor in_data(453) xor in_data(455) xor in_data(456) xor in_data(460) xor in_data(463) xor in_data(464) xor in_data(467) xor in_data(468) xor in_data(469) xor in_data(471) xor in_data(472) xor in_data(473) xor in_data(474) xor in_data(476) xor in_data(478) xor in_data(479) xor in_data(481) xor in_data(482) xor in_data(484) xor in_data(485) xor in_data(486) xor in_data(488) xor in_data(490) xor in_data(492) xor in_data(493) xor in_data(495) xor in_data(498) xor in_data(500) xor in_data(501) xor in_data(502) xor in_data(504) xor in_data(508);

out_data(23)<= in_data(5) xor in_data(8) xor in_data(10) xor in_data(15) xor in_data(16) xor in_data(17) xor in_data(18) xor in_data(21) xor in_data(24) xor in_data(25) xor in_data(27) xor in_data(28) xor in_data(29) xor in_data(33) xor in_data(34) xor in_data(35) xor in_data(38) xor in_data(42) xor in_data(45) xor in_data(50) xor in_data(53) xor in_data(54) xor in_data(55) xor in_data(57) xor in_data(59) xor in_data(60) xor in_data(61) xor in_data(62) xor in_data(63) xor in_data(64) xor in_data(65) xor in_data(67) xor in_data(69) xor in_data(72) xor in_data(76) xor in_data(77) xor in_data(79) xor in_data(80) xor in_data(82) xor in_data(84) xor in_data(90) xor in_data(91) xor in_data(94) xor in_data(95) xor in_data(98) xor in_data(100) xor in_data(103) xor in_data(105) xor in_data(107) xor in_data(111) xor in_data(113) xor in_data(116) xor in_data(117) xor in_data(118) xor in_data(122) xor in_data(124) xor in_data(126) xor in_data(127) xor in_data(128) xor in_data(131) xor in_data(133) xor in_data(135) xor in_data(136) xor in_data(144) xor in_data(145) xor in_data(147) xor in_data(148) xor in_data(149) xor in_data(150) xor in_data(154) xor in_data(158) xor in_data(160) xor in_data(161) xor in_data(163) xor in_data(165) xor in_data(166) xor in_data(169) xor in_data(172) xor in_data(175) xor in_data(177) xor in_data(178) xor in_data(181) xor in_data(182) xor in_data(184) xor in_data(185) xor in_data(189) xor in_data(190) xor in_data(192) xor in_data(195) xor in_data(196) xor in_data(197) xor in_data(198) xor in_data(205) xor in_data(206) xor in_data(207) xor in_data(208) xor in_data(209) xor in_data(211) xor in_data(212) xor in_data(215) xor in_data(217) xor in_data(218) xor in_data(220) xor in_data(221) xor in_data(222) xor in_data(223) xor in_data(224) xor in_data(229) xor in_data(231) xor in_data(233) xor in_data(235) xor in_data(237) xor in_data(238) xor in_data(239) xor in_data(240) xor in_data(242) xor in_data(243) xor in_data(244) xor in_data(245) xor in_data(246) xor in_data(247) xor in_data(250) xor in_data(251) xor in_data(252) xor in_data(253) xor in_data(255) xor in_data(258) xor in_data(261) xor in_data(262) xor in_data(263) xor in_data(264) xor in_data(265) xor in_data(268) xor in_data(270) xor in_data(271) xor in_data(272) xor in_data(273) xor in_data(274) xor in_data(276) xor in_data(283) xor in_data(285) xor in_data(286) xor in_data(290) xor in_data(293) xor in_data(294) xor in_data(297) xor in_data(298) xor in_data(299) xor in_data(301) xor in_data(302) xor in_data(303) xor in_data(304) xor in_data(306) xor in_data(308) xor in_data(309) xor in_data(311) xor in_data(312) xor in_data(314) xor in_data(315) xor in_data(316) xor in_data(318) xor in_data(320) xor in_data(322) xor in_data(323) xor in_data(325) xor in_data(328) xor in_data(330) xor in_data(331) xor in_data(332) xor in_data(334) xor in_data(338) xor in_data(344) xor in_data(349) xor in_data(350) xor in_data(352) xor in_data(354) xor in_data(355) xor in_data(356) xor in_data(358) xor in_data(359) xor in_data(364) xor in_data(368) xor in_data(369) xor in_data(370) xor in_data(371) xor in_data(372) xor in_data(373) xor in_data(374) xor in_data(375) xor in_data(376) xor in_data(380) xor in_data(381) xor in_data(387) xor in_data(389) xor in_data(393) xor in_data(394) xor in_data(395) xor in_data(397) xor in_data(398) xor in_data(400) xor in_data(405) xor in_data(407) xor in_data(408) xor in_data(409) xor in_data(414) xor in_data(415) xor in_data(416) xor in_data(422) xor in_data(423) xor in_data(424) xor in_data(426) xor in_data(429) xor in_data(430) xor in_data(432) xor in_data(434) xor in_data(436) xor in_data(439) xor in_data(440) xor in_data(444) xor in_data(445) xor in_data(446) xor in_data(447) xor in_data(449) xor in_data(450) xor in_data(452) xor in_data(453) xor in_data(456) xor in_data(457) xor in_data(458) xor in_data(459) xor in_data(460) xor in_data(461) xor in_data(463) xor in_data(464) xor in_data(465) xor in_data(467) xor in_data(468) xor in_data(469) xor in_data(472) xor in_data(473) xor in_data(474) xor in_data(477) xor in_data(478) xor in_data(483) xor in_data(484) xor in_data(488) xor in_data(490) xor in_data(491) xor in_data(492) xor in_data(493) xor in_data(496) xor in_data(497) xor in_data(499) xor in_data(503) xor in_data(504) xor in_data(507);

out_data(24)<= in_data(2) xor in_data(5) xor in_data(7) xor in_data(8) xor in_data(11) xor in_data(12) xor in_data(14) xor in_data(15) xor in_data(19) xor in_data(20) xor in_data(22) xor in_data(25) xor in_data(26) xor in_data(27) xor in_data(28) xor in_data(35) xor in_data(36) xor in_data(37) xor in_data(38) xor in_data(39) xor in_data(41) xor in_data(42) xor in_data(45) xor in_data(47) xor in_data(48) xor in_data(50) xor in_data(51) xor in_data(52) xor in_data(53) xor in_data(54) xor in_data(59) xor in_data(61) xor in_data(63) xor in_data(65) xor in_data(67) xor in_data(68) xor in_data(69) xor in_data(70) xor in_data(72) xor in_data(73) xor in_data(74) xor in_data(75) xor in_data(76) xor in_data(77) xor in_data(80) xor in_data(81) xor in_data(82) xor in_data(83) xor in_data(85) xor in_data(88) xor in_data(91) xor in_data(92) xor in_data(93) xor in_data(94) xor in_data(95) xor in_data(98) xor in_data(100) xor in_data(101) xor in_data(102) xor in_data(103) xor in_data(104) xor in_data(106) xor in_data(113) xor in_data(115) xor in_data(116) xor in_data(120) xor in_data(123) xor in_data(124) xor in_data(127) xor in_data(128) xor in_data(129) xor in_data(131) xor in_data(132) xor in_data(133) xor in_data(134) xor in_data(136) xor in_data(138) xor in_data(139) xor in_data(141) xor in_data(142) xor in_data(144) xor in_data(145) xor in_data(146) xor in_data(148) xor in_data(150) xor in_data(152) xor in_data(153) xor in_data(155) xor in_data(158) xor in_data(160) xor in_data(161) xor in_data(162) xor in_data(164) xor in_data(168) xor in_data(174) xor in_data(179) xor in_data(180) xor in_data(182) xor in_data(184) xor in_data(185) xor in_data(186) xor in_data(188) xor in_data(189) xor in_data(194) xor in_data(198) xor in_data(199) xor in_data(200) xor in_data(201) xor in_data(202) xor in_data(203) xor in_data(204) xor in_data(205) xor in_data(206) xor in_data(210) xor in_data(211) xor in_data(217) xor in_data(219) xor in_data(223) xor in_data(224) xor in_data(225) xor in_data(227) xor in_data(228) xor in_data(230) xor in_data(235) xor in_data(237) xor in_data(238) xor in_data(239) xor in_data(244) xor in_data(245) xor in_data(246) xor in_data(252) xor in_data(253) xor in_data(254) xor in_data(256) xor in_data(259) xor in_data(260) xor in_data(262) xor in_data(264) xor in_data(266) xor in_data(269) xor in_data(270) xor in_data(274) xor in_data(275) xor in_data(276) xor in_data(277) xor in_data(279) xor in_data(280) xor in_data(282) xor in_data(283) xor in_data(286) xor in_data(287) xor in_data(288) xor in_data(289) xor in_data(290) xor in_data(291) xor in_data(293) xor in_data(294) xor in_data(295) xor in_data(297) xor in_data(298) xor in_data(299) xor in_data(302) xor in_data(303) xor in_data(304) xor in_data(307) xor in_data(308) xor in_data(313) xor in_data(314) xor in_data(318) xor in_data(320) xor in_data(321) xor in_data(322) xor in_data(323) xor in_data(326) xor in_data(327) xor in_data(329) xor in_data(333) xor in_data(334) xor in_data(337) xor in_data(346) xor in_data(349) xor in_data(351) xor in_data(356) xor in_data(357) xor in_data(358) xor in_data(359) xor in_data(362) xor in_data(365) xor in_data(366) xor in_data(368) xor in_data(369) xor in_data(370) xor in_data(374) xor in_data(375) xor in_data(376) xor in_data(379) xor in_data(383) xor in_data(386) xor in_data(391) xor in_data(394) xor in_data(395) xor in_data(396) xor in_data(398) xor in_data(400) xor in_data(401) xor in_data(402) xor in_data(403) xor in_data(404) xor in_data(405) xor in_data(406) xor in_data(408) xor in_data(410) xor in_data(413) xor in_data(417) xor in_data(418) xor in_data(420) xor in_data(421) xor in_data(423) xor in_data(425) xor in_data(431) xor in_data(432) xor in_data(435) xor in_data(436) xor in_data(439) xor in_data(441) xor in_data(444) xor in_data(446) xor in_data(448) xor in_data(452) xor in_data(454) xor in_data(457) xor in_data(458) xor in_data(459) xor in_data(463) xor in_data(465) xor in_data(467) xor in_data(468) xor in_data(469) xor in_data(472) xor in_data(474) xor in_data(476) xor in_data(477) xor in_data(485) xor in_data(486) xor in_data(488) xor in_data(489) xor in_data(490) xor in_data(491) xor in_data(495) xor in_data(499) xor in_data(501) xor in_data(502) xor in_data(504) xor in_data(506) xor in_data(507) xor in_data(510);

out_data(25)<= in_data(4) xor in_data(9) xor in_data(10) xor in_data(12) xor in_data(14) xor in_data(15) xor in_data(16) xor in_data(18) xor in_data(19) xor in_data(24) xor in_data(28) xor in_data(29) xor in_data(30) xor in_data(31) xor in_data(32) xor in_data(33) xor in_data(34) xor in_data(35) xor in_data(36) xor in_data(40) xor in_data(41) xor in_data(47) xor in_data(49) xor in_data(53) xor in_data(54) xor in_data(55) xor in_data(57) xor in_data(58) xor in_data(60) xor in_data(65) xor in_data(67) xor in_data(68) xor in_data(69) xor in_data(74) xor in_data(75) xor in_data(76) xor in_data(82) xor in_data(83) xor in_data(84) xor in_data(86) xor in_data(89) xor in_data(90) xor in_data(92) xor in_data(94) xor in_data(96) xor in_data(99) xor in_data(100) xor in_data(104) xor in_data(105) xor in_data(106) xor in_data(107) xor in_data(109) xor in_data(110) xor in_data(112) xor in_data(113) xor in_data(116) xor in_data(117) xor in_data(118) xor in_data(119) xor in_data(120) xor in_data(121) xor in_data(123) xor in_data(124) xor in_data(125) xor in_data(127) xor in_data(128) xor in_data(129) xor in_data(132) xor in_data(133) xor in_data(134) xor in_data(137) xor in_data(138) xor in_data(143) xor in_data(144) xor in_data(148) xor in_data(150) xor in_data(151) xor in_data(152) xor in_data(153) xor in_data(156) xor in_data(157) xor in_data(159) xor in_data(163) xor in_data(164) xor in_data(167) xor in_data(176) xor in_data(179) xor in_data(181) xor in_data(186) xor in_data(187) xor in_data(188) xor in_data(189) xor in_data(192) xor in_data(195) xor in_data(196) xor in_data(198) xor in_data(199) xor in_data(200) xor in_data(204) xor in_data(205) xor in_data(206) xor in_data(209) xor in_data(213) xor in_data(216) xor in_data(221) xor in_data(224) xor in_data(225) xor in_data(226) xor in_data(228) xor in_data(230) xor in_data(231) xor in_data(232) xor in_data(233) xor in_data(234) xor in_data(235) xor in_data(236) xor in_data(238) xor in_data(240) xor in_data(243) xor in_data(247) xor in_data(248) xor in_data(250) xor in_data(251) xor in_data(253) xor in_data(255) xor in_data(261) xor in_data(262) xor in_data(265) xor in_data(266) xor in_data(269) xor in_data(271) xor in_data(274) xor in_data(276) xor in_data(278) xor in_data(282) xor in_data(284) xor in_data(287) xor in_data(288) xor in_data(289) xor in_data(293) xor in_data(295) xor in_data(297) xor in_data(298) xor in_data(299) xor in_data(302) xor in_data(304) xor in_data(306) xor in_data(307) xor in_data(315) xor in_data(316) xor in_data(318) xor in_data(319) xor in_data(320) xor in_data(321) xor in_data(325) xor in_data(329) xor in_data(331) xor in_data(332) xor in_data(334) xor in_data(336) xor in_data(337) xor in_data(340) xor in_data(343) xor in_data(346) xor in_data(348) xor in_data(349) xor in_data(352) xor in_data(353) xor in_data(355) xor in_data(356) xor in_data(360) xor in_data(361) xor in_data(363) xor in_data(366) xor in_data(367) xor in_data(368) xor in_data(369) xor in_data(376) xor in_data(377) xor in_data(378) xor in_data(379) xor in_data(380) xor in_data(382) xor in_data(383) xor in_data(386) xor in_data(388) xor in_data(389) xor in_data(391) xor in_data(392) xor in_data(393) xor in_data(394) xor in_data(395) xor in_data(400) xor in_data(402) xor in_data(404) xor in_data(406) xor in_data(408) xor in_data(409) xor in_data(410) xor in_data(411) xor in_data(413) xor in_data(414) xor in_data(415) xor in_data(416) xor in_data(417) xor in_data(418) xor in_data(421) xor in_data(422) xor in_data(423) xor in_data(424) xor in_data(426) xor in_data(429) xor in_data(432) xor in_data(433) xor in_data(434) xor in_data(435) xor in_data(436) xor in_data(439) xor in_data(441) xor in_data(442) xor in_data(443) xor in_data(444) xor in_data(445) xor in_data(447) xor in_data(454) xor in_data(456) xor in_data(457) xor in_data(461) xor in_data(464) xor in_data(465) xor in_data(468) xor in_data(469) xor in_data(470) xor in_data(472) xor in_data(473) xor in_data(474) xor in_data(475) xor in_data(477) xor in_data(479) xor in_data(480) xor in_data(482) xor in_data(483) xor in_data(485) xor in_data(486) xor in_data(487) xor in_data(489) xor in_data(491) xor in_data(493) xor in_data(494) xor in_data(496) xor in_data(499) xor in_data(501) xor in_data(502) xor in_data(503) xor in_data(505) xor in_data(509);

out_data(26)<= in_data(6) xor in_data(9) xor in_data(11) xor in_data(16) xor in_data(17) xor in_data(18) xor in_data(19) xor in_data(22) xor in_data(25) xor in_data(26) xor in_data(28) xor in_data(29) xor in_data(30) xor in_data(34) xor in_data(35) xor in_data(36) xor in_data(39) xor in_data(43) xor in_data(46) xor in_data(51) xor in_data(54) xor in_data(55) xor in_data(56) xor in_data(58) xor in_data(60) xor in_data(61) xor in_data(62) xor in_data(63) xor in_data(64) xor in_data(65) xor in_data(66) xor in_data(68) xor in_data(70) xor in_data(73) xor in_data(77) xor in_data(78) xor in_data(80) xor in_data(81) xor in_data(83) xor in_data(85) xor in_data(91) xor in_data(92) xor in_data(95) xor in_data(96) xor in_data(99) xor in_data(101) xor in_data(104) xor in_data(106) xor in_data(108) xor in_data(112) xor in_data(114) xor in_data(117) xor in_data(118) xor in_data(119) xor in_data(123) xor in_data(125) xor in_data(127) xor in_data(128) xor in_data(129) xor in_data(132) xor in_data(134) xor in_data(136) xor in_data(137) xor in_data(145) xor in_data(146) xor in_data(148) xor in_data(149) xor in_data(150) xor in_data(151) xor in_data(155) xor in_data(159) xor in_data(161) xor in_data(162) xor in_data(164) xor in_data(166) xor in_data(167) xor in_data(170) xor in_data(173) xor in_data(176) xor in_data(178) xor in_data(179) xor in_data(182) xor in_data(183) xor in_data(185) xor in_data(186) xor in_data(190) xor in_data(191) xor in_data(193) xor in_data(196) xor in_data(197) xor in_data(198) xor in_data(199) xor in_data(206) xor in_data(207) xor in_data(208) xor in_data(209) xor in_data(210) xor in_data(212) xor in_data(213) xor in_data(216) xor in_data(218) xor in_data(219) xor in_data(221) xor in_data(222) xor in_data(223) xor in_data(224) xor in_data(225) xor in_data(230) xor in_data(232) xor in_data(234) xor in_data(236) xor in_data(238) xor in_data(239) xor in_data(240) xor in_data(241) xor in_data(243) xor in_data(244) xor in_data(245) xor in_data(246) xor in_data(247) xor in_data(248) xor in_data(251) xor in_data(252) xor in_data(253) xor in_data(254) xor in_data(256) xor in_data(259) xor in_data(262) xor in_data(263) xor in_data(264) xor in_data(265) xor in_data(266) xor in_data(269) xor in_data(271) xor in_data(272) xor in_data(273) xor in_data(274) xor in_data(275) xor in_data(277) xor in_data(284) xor in_data(286) xor in_data(287) xor in_data(291) xor in_data(294) xor in_data(295) xor in_data(298) xor in_data(299) xor in_data(300) xor in_data(302) xor in_data(303) xor in_data(304) xor in_data(305) xor in_data(307) xor in_data(309) xor in_data(310) xor in_data(312) xor in_data(313) xor in_data(315) xor in_data(316) xor in_data(317) xor in_data(319) xor in_data(321) xor in_data(323) xor in_data(324) xor in_data(326) xor in_data(329) xor in_data(331) xor in_data(332) xor in_data(333) xor in_data(335) xor in_data(339) xor in_data(345) xor in_data(350) xor in_data(351) xor in_data(353) xor in_data(355) xor in_data(356) xor in_data(357) xor in_data(359) xor in_data(360) xor in_data(365) xor in_data(369) xor in_data(370) xor in_data(371) xor in_data(372) xor in_data(373) xor in_data(374) xor in_data(375) xor in_data(376) xor in_data(377) xor in_data(381) xor in_data(382) xor in_data(388) xor in_data(390) xor in_data(394) xor in_data(395) xor in_data(396) xor in_data(398) xor in_data(399) xor in_data(401) xor in_data(406) xor in_data(408) xor in_data(409) xor in_data(410) xor in_data(415) xor in_data(416) xor in_data(417) xor in_data(423) xor in_data(424) xor in_data(425) xor in_data(427) xor in_data(430) xor in_data(431) xor in_data(433) xor in_data(435) xor in_data(437) xor in_data(440) xor in_data(441) xor in_data(445) xor in_data(446) xor in_data(447) xor in_data(448) xor in_data(450) xor in_data(451) xor in_data(453) xor in_data(454) xor in_data(457) xor in_data(458) xor in_data(459) xor in_data(460) xor in_data(461) xor in_data(462) xor in_data(464) xor in_data(465) xor in_data(466) xor in_data(468) xor in_data(469) xor in_data(470) xor in_data(473) xor in_data(474) xor in_data(475) xor in_data(478) xor in_data(479) xor in_data(484) xor in_data(485) xor in_data(489) xor in_data(491) xor in_data(492) xor in_data(493) xor in_data(494) xor in_data(497) xor in_data(498) xor in_data(500) xor in_data(504) xor in_data(505) xor in_data(508);

out_data(27)<='0';

out_data(28)<='0';

out_data(29)<='0';

out_data(30)<='0';

out_data(31)<='0';

out_data(32)<='0';

out_data(33)<='0';

out_data(34)<='0';

out_data(35)<='0';

out_data(36)<= in_data(0) xor in_data(9) xor in_data(10) xor in_data(11) xor in_data(12) xor in_data(17) xor in_data(19) xor in_data(22) xor in_data(24) xor in_data(25) xor in_data(26) xor in_data(33) xor in_data(35) xor in_data(36) xor in_data(38) xor in_data(41) xor in_data(42) xor in_data(44) xor in_data(45) xor in_data(46) xor in_data(47) xor in_data(50) xor in_data(52) xor in_data(57) xor in_data(58) xor in_data(63) xor in_data(64) xor in_data(65) xor in_data(70) xor in_data(71) xor in_data(73) xor in_data(74) xor in_data(75) xor in_data(77) xor in_data(78) xor in_data(81) xor in_data(84) xor in_data(87) xor in_data(89) xor in_data(91) xor in_data(94) xor in_data(99) xor in_data(104) xor in_data(105) xor in_data(106) xor in_data(107) xor in_data(108) xor in_data(109) xor in_data(110) xor in_data(111) xor in_data(112) xor in_data(114) xor in_data(116) xor in_data(117) xor in_data(118) xor in_data(119) xor in_data(120) xor in_data(123) xor in_data(124) xor in_data(125) xor in_data(128) xor in_data(130) xor in_data(131) xor in_data(132) xor in_data(133) xor in_data(134) xor in_data(135) xor in_data(136) xor in_data(139) xor in_data(142) xor in_data(143) xor in_data(144) xor in_data(146) xor in_data(147) xor in_data(149) xor in_data(151) xor in_data(152) xor in_data(153) xor in_data(156) xor in_data(157) xor in_data(158) xor in_data(159) xor in_data(160) xor in_data(162) xor in_data(163) xor in_data(164) xor in_data(165) xor in_data(166) xor in_data(168) xor in_data(174) xor in_data(177) xor in_data(179) xor in_data(180) xor in_data(182) xor in_data(183) xor in_data(184) xor in_data(188) xor in_data(189) xor in_data(190) xor in_data(193) xor in_data(194) xor in_data(198) xor in_data(199) xor in_data(200) xor in_data(201) xor in_data(202) xor in_data(208) xor in_data(210) xor in_data(212) xor in_data(214) xor in_data(216) xor in_data(217) xor in_data(220) xor in_data(222) xor in_data(224) xor in_data(225) xor in_data(226) xor in_data(228) xor in_data(232) xor in_data(233) xor in_data(235) xor in_data(237) xor in_data(239) xor in_data(243) xor in_data(244) xor in_data(245) xor in_data(247) xor in_data(250) xor in_data(253) xor in_data(254) xor in_data(256) xor in_data(260) xor in_data(262) xor in_data(264) xor in_data(265) xor in_data(267) xor in_data(269) xor in_data(272) xor in_data(273) xor in_data(274) xor in_data(275) xor in_data(276) xor in_data(277) xor in_data(281) xor in_data(282) xor in_data(284) xor in_data(285) xor in_data(287) xor in_data(292) xor in_data(294) xor in_data(295) xor in_data(296) xor in_data(298) xor in_data(299) xor in_data(300) xor in_data(301) xor in_data(303) xor in_data(305) xor in_data(312) xor in_data(313) xor in_data(316) xor in_data(317) xor in_data(320) xor in_data(324) xor in_data(325) xor in_data(328) xor in_data(330) xor in_data(331) xor in_data(336) xor in_data(339) xor in_data(340) xor in_data(343) xor in_data(344) xor in_data(345) xor in_data(346) xor in_data(348) xor in_data(351) xor in_data(352) xor in_data(353) xor in_data(357) xor in_data(360) xor in_data(361) xor in_data(362) xor in_data(363) xor in_data(366) xor in_data(367) xor in_data(369) xor in_data(370) xor in_data(373) xor in_data(374) xor in_data(375) xor in_data(377) xor in_data(379) xor in_data(381) xor in_data(382) xor in_data(383) xor in_data(384) xor in_data(386) xor in_data(387) xor in_data(389) xor in_data(390) xor in_data(396) xor in_data(397) xor in_data(399) xor in_data(402) xor in_data(404) xor in_data(407) xor in_data(408) xor in_data(416) xor in_data(420) xor in_data(424) xor in_data(425) xor in_data(426) xor in_data(427) xor in_data(429) xor in_data(430) xor in_data(431) xor in_data(434) xor in_data(440) xor in_data(441) xor in_data(442) xor in_data(444) xor in_data(445) xor in_data(446) xor in_data(448) xor in_data(450) xor in_data(451) xor in_data(455) xor in_data(457) xor in_data(458) xor in_data(459) xor in_data(460) xor in_data(464) xor in_data(466) xor in_data(470) xor in_data(473) xor in_data(477) xor in_data(479) xor in_data(480) xor in_data(483) xor in_data(484) xor in_data(486) xor in_data(488) xor in_data(489) xor in_data(491) xor in_data(492) xor in_data(494) xor in_data(495) xor in_data(496) xor in_data(497) xor in_data(498) xor in_data(499) xor in_data(501) xor in_data(502) xor in_data(506) xor in_data(507);

out_data(37)<= in_data(2) xor in_data(3) xor in_data(4) xor in_data(5) xor in_data(6) xor in_data(7) xor in_data(8) xor in_data(9) xor in_data(10) xor in_data(12) xor in_data(14) xor in_data(15) xor in_data(16) xor in_data(17) xor in_data(18) xor in_data(21) xor in_data(22) xor in_data(23) xor in_data(26) xor in_data(28) xor in_data(29) xor in_data(30) xor in_data(31) xor in_data(32) xor in_data(33) xor in_data(34) xor in_data(37) xor in_data(40) xor in_data(41) xor in_data(42) xor in_data(44) xor in_data(45) xor in_data(47) xor in_data(49) xor in_data(50) xor in_data(51) xor in_data(54) xor in_data(55) xor in_data(56) xor in_data(57) xor in_data(58) xor in_data(60) xor in_data(61) xor in_data(62) xor in_data(63) xor in_data(64) xor in_data(66) xor in_data(72) xor in_data(75) xor in_data(77) xor in_data(78) xor in_data(80) xor in_data(81) xor in_data(82) xor in_data(86) xor in_data(87) xor in_data(88) xor in_data(91) xor in_data(92) xor in_data(96) xor in_data(97) xor in_data(98) xor in_data(99) xor in_data(100) xor in_data(106) xor in_data(108) xor in_data(110) xor in_data(112) xor in_data(114) xor in_data(115) xor in_data(118) xor in_data(120) xor in_data(122) xor in_data(123) xor in_data(124) xor in_data(126) xor in_data(130) xor in_data(131) xor in_data(133) xor in_data(135) xor in_data(137) xor in_data(141) xor in_data(142) xor in_data(143) xor in_data(145) xor in_data(148) xor in_data(151) xor in_data(152) xor in_data(154) xor in_data(158) xor in_data(160) xor in_data(162) xor in_data(163) xor in_data(165) xor in_data(167) xor in_data(170) xor in_data(171) xor in_data(172) xor in_data(173) xor in_data(174) xor in_data(175) xor in_data(179) xor in_data(180) xor in_data(182) xor in_data(183) xor in_data(185) xor in_data(190) xor in_data(192) xor in_data(193) xor in_data(194) xor in_data(196) xor in_data(197) xor in_data(198) xor in_data(199) xor in_data(201) xor in_data(203) xor in_data(210) xor in_data(211) xor in_data(214) xor in_data(215) xor in_data(218) xor in_data(222) xor in_data(223) xor in_data(226) xor in_data(228) xor in_data(229) xor in_data(234) xor in_data(237) xor in_data(238) xor in_data(241) xor in_data(242) xor in_data(243) xor in_data(244) xor in_data(246) xor in_data(249) xor in_data(250) xor in_data(251) xor in_data(255) xor in_data(258) xor in_data(259) xor in_data(260) xor in_data(261) xor in_data(264) xor in_data(265) xor in_data(267) xor in_data(268) xor in_data(271) xor in_data(272) xor in_data(273) xor in_data(275) xor in_data(277) xor in_data(279) xor in_data(280) xor in_data(281) xor in_data(282) xor in_data(284) xor in_data(285) xor in_data(287) xor in_data(288) xor in_data(294) xor in_data(295) xor in_data(297) xor in_data(300) xor in_data(302) xor in_data(305) xor in_data(306) xor in_data(314) xor in_data(318) xor in_data(322) xor in_data(323) xor in_data(324) xor in_data(325) xor in_data(327) xor in_data(328) xor in_data(329) xor in_data(332) xor in_data(338) xor in_data(339) xor in_data(340) xor in_data(342) xor in_data(343) xor in_data(344) xor in_data(346) xor in_data(348) xor in_data(349) xor in_data(353) xor in_data(355) xor in_data(356) xor in_data(357) xor in_data(358) xor in_data(362) xor in_data(364) xor in_data(368) xor in_data(371) xor in_data(375) xor in_data(377) xor in_data(378) xor in_data(381) xor in_data(382) xor in_data(384) xor in_data(386) xor in_data(387) xor in_data(389) xor in_data(390) xor in_data(392) xor in_data(393) xor in_data(394) xor in_data(395) xor in_data(396) xor in_data(397) xor in_data(399) xor in_data(400) xor in_data(404) xor in_data(405) xor in_data(409) xor in_data(418) xor in_data(419) xor in_data(420) xor in_data(421) xor in_data(426) xor in_data(428) xor in_data(431) xor in_data(433) xor in_data(434) xor in_data(435) xor in_data(442) xor in_data(444) xor in_data(445) xor in_data(447) xor in_data(450) xor in_data(451) xor in_data(453) xor in_data(454) xor in_data(455) xor in_data(456) xor in_data(459) xor in_data(461) xor in_data(466) xor in_data(467) xor in_data(472) xor in_data(473) xor in_data(474) xor in_data(479) xor in_data(480) xor in_data(482) xor in_data(483) xor in_data(484) xor in_data(486) xor in_data(487) xor in_data(490) xor in_data(493) xor in_data(496) xor in_data(498) xor in_data(500) xor in_data(503) xor in_data(508);

out_data(38)<= in_data(4) xor in_data(6) xor in_data(8) xor in_data(10) xor in_data(12) xor in_data(13) xor in_data(16) xor in_data(18) xor in_data(20) xor in_data(21) xor in_data(22) xor in_data(24) xor in_data(28) xor in_data(29) xor in_data(31) xor in_data(33) xor in_data(35) xor in_data(39) xor in_data(40) xor in_data(41) xor in_data(43) xor in_data(46) xor in_data(49) xor in_data(50) xor in_data(52) xor in_data(56) xor in_data(58) xor in_data(60) xor in_data(61) xor in_data(63) xor in_data(65) xor in_data(68) xor in_data(69) xor in_data(70) xor in_data(71) xor in_data(72) xor in_data(73) xor in_data(77) xor in_data(78) xor in_data(80) xor in_data(81) xor in_data(83) xor in_data(88) xor in_data(90) xor in_data(91) xor in_data(92) xor in_data(94) xor in_data(95) xor in_data(96) xor in_data(97) xor in_data(99) xor in_data(101) xor in_data(108) xor in_data(109) xor in_data(112) xor in_data(113) xor in_data(116) xor in_data(120) xor in_data(121) xor in_data(124) xor in_data(126) xor in_data(127) xor in_data(132) xor in_data(135) xor in_data(136) xor in_data(139) xor in_data(140) xor in_data(141) xor in_data(142) xor in_data(144) xor in_data(147) xor in_data(148) xor in_data(149) xor in_data(153) xor in_data(156) xor in_data(157) xor in_data(158) xor in_data(159) xor in_data(162) xor in_data(163) xor in_data(165) xor in_data(166) xor in_data(169) xor in_data(170) xor in_data(171) xor in_data(173) xor in_data(175) xor in_data(177) xor in_data(178) xor in_data(179) xor in_data(180) xor in_data(182) xor in_data(183) xor in_data(185) xor in_data(186) xor in_data(192) xor in_data(193) xor in_data(195) xor in_data(198) xor in_data(200) xor in_data(203) xor in_data(204) xor in_data(212) xor in_data(216) xor in_data(220) xor in_data(221) xor in_data(222) xor in_data(223) xor in_data(225) xor in_data(226) xor in_data(227) xor in_data(230) xor in_data(236) xor in_data(237) xor in_data(238) xor in_data(240) xor in_data(241) xor in_data(242) xor in_data(244) xor in_data(246) xor in_data(247) xor in_data(251) xor in_data(253) xor in_data(254) xor in_data(255) xor in_data(256) xor in_data(260) xor in_data(262) xor in_data(266) xor in_data(269) xor in_data(273) xor in_data(275) xor in_data(276) xor in_data(279) xor in_data(280) xor in_data(282) xor in_data(284) xor in_data(285) xor in_data(287) xor in_data(288) xor in_data(290) xor in_data(291) xor in_data(292) xor in_data(293) xor in_data(294) xor in_data(295) xor in_data(297) xor in_data(298) xor in_data(302) xor in_data(303) xor in_data(307) xor in_data(316) xor in_data(317) xor in_data(318) xor in_data(319) xor in_data(324) xor in_data(326) xor in_data(329) xor in_data(331) xor in_data(332) xor in_data(333) xor in_data(340) xor in_data(342) xor in_data(343) xor in_data(345) xor in_data(348) xor in_data(349) xor in_data(351) xor in_data(352) xor in_data(353) xor in_data(354) xor in_data(357) xor in_data(359) xor in_data(364) xor in_data(365) xor in_data(370) xor in_data(371) xor in_data(372) xor in_data(377) xor in_data(378) xor in_data(380) xor in_data(381) xor in_data(382) xor in_data(384) xor in_data(385) xor in_data(388) xor in_data(391) xor in_data(394) xor in_data(396) xor in_data(398) xor in_data(401) xor in_data(406) xor in_data(411) xor in_data(412) xor in_data(413) xor in_data(414) xor in_data(415) xor in_data(416) xor in_data(417) xor in_data(418) xor in_data(419) xor in_data(421) xor in_data(423) xor in_data(424) xor in_data(425) xor in_data(426) xor in_data(427) xor in_data(430) xor in_data(431) xor in_data(432) xor in_data(435) xor in_data(437) xor in_data(438) xor in_data(439) xor in_data(440) xor in_data(441) xor in_data(442) xor in_data(443) xor in_data(446) xor in_data(449) xor in_data(450) xor in_data(451) xor in_data(453) xor in_data(454) xor in_data(456) xor in_data(458) xor in_data(459) xor in_data(460) xor in_data(463) xor in_data(464) xor in_data(465) xor in_data(466) xor in_data(467) xor in_data(469) xor in_data(470) xor in_data(471) xor in_data(472) xor in_data(473) xor in_data(475) xor in_data(481) xor in_data(484) xor in_data(486) xor in_data(487) xor in_data(489) xor in_data(490) xor in_data(491) xor in_data(495) xor in_data(496) xor in_data(497) xor in_data(500) xor in_data(501) xor in_data(505) xor in_data(506) xor in_data(507) xor in_data(508) xor in_data(509);

out_data(39)<= in_data(6) xor in_data(7) xor in_data(10) xor in_data(11) xor in_data(14) xor in_data(18) xor in_data(19) xor in_data(22) xor in_data(24) xor in_data(25) xor in_data(30) xor in_data(33) xor in_data(34) xor in_data(37) xor in_data(38) xor in_data(39) xor in_data(40) xor in_data(42) xor in_data(45) xor in_data(46) xor in_data(47) xor in_data(51) xor in_data(54) xor in_data(55) xor in_data(56) xor in_data(57) xor in_data(60) xor in_data(61) xor in_data(63) xor in_data(64) xor in_data(67) xor in_data(68) xor in_data(69) xor in_data(71) xor in_data(73) xor in_data(75) xor in_data(76) xor in_data(77) xor in_data(78) xor in_data(80) xor in_data(81) xor in_data(83) xor in_data(84) xor in_data(90) xor in_data(91) xor in_data(93) xor in_data(96) xor in_data(98) xor in_data(101) xor in_data(102) xor in_data(110) xor in_data(114) xor in_data(118) xor in_data(119) xor in_data(120) xor in_data(121) xor in_data(123) xor in_data(124) xor in_data(125) xor in_data(128) xor in_data(134) xor in_data(135) xor in_data(136) xor in_data(138) xor in_data(139) xor in_data(140) xor in_data(142) xor in_data(144) xor in_data(145) xor in_data(149) xor in_data(151) xor in_data(152) xor in_data(153) xor in_data(154) xor in_data(158) xor in_data(160) xor in_data(164) xor in_data(167) xor in_data(171) xor in_data(173) xor in_data(174) xor in_data(177) xor in_data(178) xor in_data(180) xor in_data(182) xor in_data(183) xor in_data(185) xor in_data(186) xor in_data(188) xor in_data(189) xor in_data(190) xor in_data(191) xor in_data(192) xor in_data(193) xor in_data(195) xor in_data(196) xor in_data(200) xor in_data(201) xor in_data(205) xor in_data(214) xor in_data(215) xor in_data(216) xor in_data(217) xor in_data(222) xor in_data(224) xor in_data(227) xor in_data(229) xor in_data(230) xor in_data(231) xor in_data(238) xor in_data(240) xor in_data(241) xor in_data(243) xor in_data(246) xor in_data(247) xor in_data(249) xor in_data(250) xor in_data(251) xor in_data(252) xor in_data(255) xor in_data(257) xor in_data(262) xor in_data(263) xor in_data(268) xor in_data(269) xor in_data(270) xor in_data(275) xor in_data(276) xor in_data(278) xor in_data(279) xor in_data(280) xor in_data(282) xor in_data(283) xor in_data(286) xor in_data(289) xor in_data(292) xor in_data(294) xor in_data(296) xor in_data(299) xor in_data(304) xor in_data(309) xor in_data(310) xor in_data(311) xor in_data(312) xor in_data(313) xor in_data(314) xor in_data(315) xor in_data(316) xor in_data(317) xor in_data(319) xor in_data(321) xor in_data(322) xor in_data(323) xor in_data(324) xor in_data(325) xor in_data(328) xor in_data(329) xor in_data(330) xor in_data(333) xor in_data(335) xor in_data(336) xor in_data(337) xor in_data(338) xor in_data(339) xor in_data(340) xor in_data(341) xor in_data(344) xor in_data(347) xor in_data(348) xor in_data(349) xor in_data(351) xor in_data(352) xor in_data(354) xor in_data(356) xor in_data(357) xor in_data(358) xor in_data(361) xor in_data(362) xor in_data(363) xor in_data(364) xor in_data(365) xor in_data(367) xor in_data(368) xor in_data(369) xor in_data(370) xor in_data(371) xor in_data(373) xor in_data(379) xor in_data(382) xor in_data(384) xor in_data(385) xor in_data(387) xor in_data(388) xor in_data(389) xor in_data(393) xor in_data(394) xor in_data(395) xor in_data(398) xor in_data(399) xor in_data(403) xor in_data(404) xor in_data(405) xor in_data(406) xor in_data(407) xor in_data(413) xor in_data(415) xor in_data(417) xor in_data(419) xor in_data(421) xor in_data(422) xor in_data(425) xor in_data(427) xor in_data(429) xor in_data(430) xor in_data(431) xor in_data(433) xor in_data(437) xor in_data(438) xor in_data(440) xor in_data(442) xor in_data(444) xor in_data(448) xor in_data(449) xor in_data(450) xor in_data(452) xor in_data(455) xor in_data(458) xor in_data(459) xor in_data(461) xor in_data(465) xor in_data(467) xor in_data(469) xor in_data(470) xor in_data(472) xor in_data(474) xor in_data(477) xor in_data(478) xor in_data(479) xor in_data(480) xor in_data(481) xor in_data(482) xor in_data(486) xor in_data(487) xor in_data(489) xor in_data(490) xor in_data(492) xor in_data(497) xor in_data(499) xor in_data(500) xor in_data(501) xor in_data(503) xor in_data(504) xor in_data(505) xor in_data(506) xor in_data(508) xor in_data(510);

out_data(40)<= in_data(8) xor in_data(9) xor in_data(10) xor in_data(11) xor in_data(16) xor in_data(18) xor in_data(21) xor in_data(23) xor in_data(24) xor in_data(25) xor in_data(32) xor in_data(34) xor in_data(35) xor in_data(37) xor in_data(40) xor in_data(41) xor in_data(43) xor in_data(44) xor in_data(45) xor in_data(46) xor in_data(49) xor in_data(51) xor in_data(56) xor in_data(57) xor in_data(62) xor in_data(63) xor in_data(64) xor in_data(69) xor in_data(70) xor in_data(72) xor in_data(73) xor in_data(74) xor in_data(76) xor in_data(77) xor in_data(80) xor in_data(83) xor in_data(86) xor in_data(88) xor in_data(90) xor in_data(93) xor in_data(98) xor in_data(103) xor in_data(104) xor in_data(105) xor in_data(106) xor in_data(107) xor in_data(108) xor in_data(109) xor in_data(110) xor in_data(111) xor in_data(113) xor in_data(115) xor in_data(116) xor in_data(117) xor in_data(118) xor in_data(119) xor in_data(122) xor in_data(123) xor in_data(124) xor in_data(127) xor in_data(129) xor in_data(130) xor in_data(131) xor in_data(132) xor in_data(133) xor in_data(134) xor in_data(135) xor in_data(138) xor in_data(141) xor in_data(142) xor in_data(143) xor in_data(145) xor in_data(146) xor in_data(148) xor in_data(150) xor in_data(151) xor in_data(152) xor in_data(155) xor in_data(156) xor in_data(157) xor in_data(158) xor in_data(159) xor in_data(161) xor in_data(162) xor in_data(163) xor in_data(164) xor in_data(165) xor in_data(167) xor in_data(173) xor in_data(176) xor in_data(178) xor in_data(179) xor in_data(181) xor in_data(182) xor in_data(183) xor in_data(187) xor in_data(188) xor in_data(189) xor in_data(192) xor in_data(193) xor in_data(197) xor in_data(198) xor in_data(199) xor in_data(200) xor in_data(201) xor in_data(207) xor in_data(209) xor in_data(211) xor in_data(213) xor in_data(215) xor in_data(216) xor in_data(219) xor in_data(221) xor in_data(223) xor in_data(224) xor in_data(225) xor in_data(227) xor in_data(231) xor in_data(232) xor in_data(234) xor in_data(236) xor in_data(238) xor in_data(242) xor in_data(243) xor in_data(244) xor in_data(246) xor in_data(249) xor in_data(252) xor in_data(253) xor in_data(255) xor in_data(259) xor in_data(261) xor in_data(263) xor in_data(264) xor in_data(266) xor in_data(268) xor in_data(271) xor in_data(272) xor in_data(273) xor in_data(274) xor in_data(275) xor in_data(276) xor in_data(280) xor in_data(281) xor in_data(283) xor in_data(284) xor in_data(286) xor in_data(291) xor in_data(293) xor in_data(294) xor in_data(295) xor in_data(297) xor in_data(298) xor in_data(299) xor in_data(300) xor in_data(302) xor in_data(304) xor in_data(311) xor in_data(312) xor in_data(315) xor in_data(316) xor in_data(319) xor in_data(323) xor in_data(324) xor in_data(327) xor in_data(329) xor in_data(330) xor in_data(335) xor in_data(338) xor in_data(339) xor in_data(342) xor in_data(343) xor in_data(344) xor in_data(345) xor in_data(347) xor in_data(350) xor in_data(351) xor in_data(352) xor in_data(356) xor in_data(359) xor in_data(360) xor in_data(361) xor in_data(362) xor in_data(365) xor in_data(366) xor in_data(368) xor in_data(369) xor in_data(372) xor in_data(373) xor in_data(374) xor in_data(376) xor in_data(378) xor in_data(380) xor in_data(381) xor in_data(382) xor in_data(383) xor in_data(385) xor in_data(386) xor in_data(388) xor in_data(389) xor in_data(395) xor in_data(396) xor in_data(398) xor in_data(401) xor in_data(403) xor in_data(406) xor in_data(407) xor in_data(415) xor in_data(419) xor in_data(423) xor in_data(424) xor in_data(425) xor in_data(426) xor in_data(428) xor in_data(429) xor in_data(430) xor in_data(433) xor in_data(439) xor in_data(440) xor in_data(441) xor in_data(443) xor in_data(444) xor in_data(445) xor in_data(447) xor in_data(449) xor in_data(450) xor in_data(454) xor in_data(456) xor in_data(457) xor in_data(458) xor in_data(459) xor in_data(463) xor in_data(465) xor in_data(469) xor in_data(472) xor in_data(476) xor in_data(478) xor in_data(479) xor in_data(482) xor in_data(483) xor in_data(485) xor in_data(487) xor in_data(488) xor in_data(490) xor in_data(491) xor in_data(493) xor in_data(494) xor in_data(495) xor in_data(496) xor in_data(497) xor in_data(498) xor in_data(500) xor in_data(501) xor in_data(505) xor in_data(506) xor in_data(510);

out_data(41)<= in_data(1) xor in_data(2) xor in_data(3) xor in_data(4) xor in_data(5) xor in_data(6) xor in_data(7) xor in_data(8) xor in_data(9) xor in_data(11) xor in_data(13) xor in_data(14) xor in_data(15) xor in_data(16) xor in_data(17) xor in_data(20) xor in_data(21) xor in_data(22) xor in_data(25) xor in_data(27) xor in_data(28) xor in_data(29) xor in_data(30) xor in_data(31) xor in_data(32) xor in_data(33) xor in_data(36) xor in_data(39) xor in_data(40) xor in_data(41) xor in_data(43) xor in_data(44) xor in_data(46) xor in_data(48) xor in_data(49) xor in_data(50) xor in_data(53) xor in_data(54) xor in_data(55) xor in_data(56) xor in_data(57) xor in_data(59) xor in_data(60) xor in_data(61) xor in_data(62) xor in_data(63) xor in_data(65) xor in_data(71) xor in_data(74) xor in_data(76) xor in_data(77) xor in_data(79) xor in_data(80) xor in_data(81) xor in_data(85) xor in_data(86) xor in_data(87) xor in_data(90) xor in_data(91) xor in_data(95) xor in_data(96) xor in_data(97) xor in_data(98) xor in_data(99) xor in_data(105) xor in_data(107) xor in_data(109) xor in_data(111) xor in_data(113) xor in_data(114) xor in_data(117) xor in_data(119) xor in_data(121) xor in_data(122) xor in_data(123) xor in_data(125) xor in_data(129) xor in_data(130) xor in_data(132) xor in_data(134) xor in_data(136) xor in_data(140) xor in_data(141) xor in_data(142) xor in_data(144) xor in_data(147) xor in_data(150) xor in_data(151) xor in_data(153) xor in_data(157) xor in_data(159) xor in_data(161) xor in_data(162) xor in_data(164) xor in_data(166) xor in_data(169) xor in_data(170) xor in_data(171) xor in_data(172) xor in_data(173) xor in_data(174) xor in_data(178) xor in_data(179) xor in_data(181) xor in_data(182) xor in_data(184) xor in_data(189) xor in_data(191) xor in_data(192) xor in_data(193) xor in_data(195) xor in_data(196) xor in_data(197) xor in_data(198) xor in_data(200) xor in_data(202) xor in_data(209) xor in_data(210) xor in_data(213) xor in_data(214) xor in_data(217) xor in_data(221) xor in_data(222) xor in_data(225) xor in_data(227) xor in_data(228) xor in_data(233) xor in_data(236) xor in_data(237) xor in_data(240) xor in_data(241) xor in_data(242) xor in_data(243) xor in_data(245) xor in_data(248) xor in_data(249) xor in_data(250) xor in_data(254) xor in_data(257) xor in_data(258) xor in_data(259) xor in_data(260) xor in_data(263) xor in_data(264) xor in_data(266) xor in_data(267) xor in_data(270) xor in_data(271) xor in_data(272) xor in_data(274) xor in_data(276) xor in_data(278) xor in_data(279) xor in_data(280) xor in_data(281) xor in_data(283) xor in_data(284) xor in_data(286) xor in_data(287) xor in_data(293) xor in_data(294) xor in_data(296) xor in_data(299) xor in_data(301) xor in_data(304) xor in_data(305) xor in_data(313) xor in_data(317) xor in_data(321) xor in_data(322) xor in_data(323) xor in_data(324) xor in_data(326) xor in_data(327) xor in_data(328) xor in_data(331) xor in_data(337) xor in_data(338) xor in_data(339) xor in_data(341) xor in_data(342) xor in_data(343) xor in_data(345) xor in_data(347) xor in_data(348) xor in_data(352) xor in_data(354) xor in_data(355) xor in_data(356) xor in_data(357) xor in_data(361) xor in_data(363) xor in_data(367) xor in_data(370) xor in_data(374) xor in_data(376) xor in_data(377) xor in_data(380) xor in_data(381) xor in_data(383) xor in_data(385) xor in_data(386) xor in_data(388) xor in_data(389) xor in_data(391) xor in_data(392) xor in_data(393) xor in_data(394) xor in_data(395) xor in_data(396) xor in_data(398) xor in_data(399) xor in_data(403) xor in_data(404) xor in_data(408) xor in_data(417) xor in_data(418) xor in_data(419) xor in_data(420) xor in_data(425) xor in_data(427) xor in_data(430) xor in_data(432) xor in_data(433) xor in_data(434) xor in_data(441) xor in_data(443) xor in_data(444) xor in_data(446) xor in_data(449) xor in_data(450) xor in_data(452) xor in_data(453) xor in_data(454) xor in_data(455) xor in_data(458) xor in_data(460) xor in_data(465) xor in_data(466) xor in_data(471) xor in_data(472) xor in_data(473) xor in_data(478) xor in_data(479) xor in_data(481) xor in_data(482) xor in_data(483) xor in_data(485) xor in_data(486) xor in_data(489) xor in_data(492) xor in_data(495) xor in_data(497) xor in_data(499) xor in_data(502) xor in_data(507);

out_data(42)<= in_data(3) xor in_data(5) xor in_data(7) xor in_data(9) xor in_data(11) xor in_data(12) xor in_data(15) xor in_data(17) xor in_data(19) xor in_data(20) xor in_data(21) xor in_data(23) xor in_data(27) xor in_data(28) xor in_data(30) xor in_data(32) xor in_data(34) xor in_data(38) xor in_data(39) xor in_data(40) xor in_data(42) xor in_data(45) xor in_data(48) xor in_data(49) xor in_data(51) xor in_data(55) xor in_data(57) xor in_data(59) xor in_data(60) xor in_data(62) xor in_data(64) xor in_data(67) xor in_data(68) xor in_data(69) xor in_data(70) xor in_data(71) xor in_data(72) xor in_data(76) xor in_data(77) xor in_data(79) xor in_data(80) xor in_data(82) xor in_data(87) xor in_data(89) xor in_data(90) xor in_data(91) xor in_data(93) xor in_data(94) xor in_data(95) xor in_data(96) xor in_data(98) xor in_data(100) xor in_data(107) xor in_data(108) xor in_data(111) xor in_data(112) xor in_data(115) xor in_data(119) xor in_data(120) xor in_data(123) xor in_data(125) xor in_data(126) xor in_data(131) xor in_data(134) xor in_data(135) xor in_data(138) xor in_data(139) xor in_data(140) xor in_data(141) xor in_data(143) xor in_data(146) xor in_data(147) xor in_data(148) xor in_data(152) xor in_data(155) xor in_data(156) xor in_data(157) xor in_data(158) xor in_data(161) xor in_data(162) xor in_data(164) xor in_data(165) xor in_data(168) xor in_data(169) xor in_data(170) xor in_data(172) xor in_data(174) xor in_data(176) xor in_data(177) xor in_data(178) xor in_data(179) xor in_data(181) xor in_data(182) xor in_data(184) xor in_data(185) xor in_data(191) xor in_data(192) xor in_data(194) xor in_data(197) xor in_data(199) xor in_data(202) xor in_data(203) xor in_data(211) xor in_data(215) xor in_data(219) xor in_data(220) xor in_data(221) xor in_data(222) xor in_data(224) xor in_data(225) xor in_data(226) xor in_data(229) xor in_data(235) xor in_data(236) xor in_data(237) xor in_data(239) xor in_data(240) xor in_data(241) xor in_data(243) xor in_data(245) xor in_data(246) xor in_data(250) xor in_data(252) xor in_data(253) xor in_data(254) xor in_data(255) xor in_data(259) xor in_data(261) xor in_data(265) xor in_data(268) xor in_data(272) xor in_data(274) xor in_data(275) xor in_data(278) xor in_data(279) xor in_data(281) xor in_data(283) xor in_data(284) xor in_data(286) xor in_data(287) xor in_data(289) xor in_data(290) xor in_data(291) xor in_data(292) xor in_data(293) xor in_data(294) xor in_data(296) xor in_data(297) xor in_data(301) xor in_data(302) xor in_data(306) xor in_data(315) xor in_data(316) xor in_data(317) xor in_data(318) xor in_data(323) xor in_data(325) xor in_data(328) xor in_data(330) xor in_data(331) xor in_data(332) xor in_data(339) xor in_data(341) xor in_data(342) xor in_data(344) xor in_data(347) xor in_data(348) xor in_data(350) xor in_data(351) xor in_data(352) xor in_data(353) xor in_data(356) xor in_data(358) xor in_data(363) xor in_data(364) xor in_data(369) xor in_data(370) xor in_data(371) xor in_data(376) xor in_data(377) xor in_data(379) xor in_data(380) xor in_data(381) xor in_data(383) xor in_data(384) xor in_data(387) xor in_data(390) xor in_data(393) xor in_data(395) xor in_data(397) xor in_data(400) xor in_data(405) xor in_data(410) xor in_data(411) xor in_data(412) xor in_data(413) xor in_data(414) xor in_data(415) xor in_data(416) xor in_data(417) xor in_data(418) xor in_data(420) xor in_data(422) xor in_data(423) xor in_data(424) xor in_data(425) xor in_data(426) xor in_data(429) xor in_data(430) xor in_data(431) xor in_data(434) xor in_data(436) xor in_data(437) xor in_data(438) xor in_data(439) xor in_data(440) xor in_data(441) xor in_data(442) xor in_data(445) xor in_data(448) xor in_data(449) xor in_data(450) xor in_data(452) xor in_data(453) xor in_data(455) xor in_data(457) xor in_data(458) xor in_data(459) xor in_data(462) xor in_data(463) xor in_data(464) xor in_data(465) xor in_data(466) xor in_data(468) xor in_data(469) xor in_data(470) xor in_data(471) xor in_data(472) xor in_data(474) xor in_data(480) xor in_data(483) xor in_data(485) xor in_data(486) xor in_data(488) xor in_data(489) xor in_data(490) xor in_data(494) xor in_data(495) xor in_data(496) xor in_data(499) xor in_data(500) xor in_data(504) xor in_data(505) xor in_data(506) xor in_data(507) xor in_data(508);

out_data(43)<= in_data(5) xor in_data(6) xor in_data(9) xor in_data(10) xor in_data(13) xor in_data(17) xor in_data(18) xor in_data(21) xor in_data(23) xor in_data(24) xor in_data(29) xor in_data(32) xor in_data(33) xor in_data(36) xor in_data(37) xor in_data(38) xor in_data(39) xor in_data(41) xor in_data(44) xor in_data(45) xor in_data(46) xor in_data(50) xor in_data(53) xor in_data(54) xor in_data(55) xor in_data(56) xor in_data(59) xor in_data(60) xor in_data(62) xor in_data(63) xor in_data(66) xor in_data(67) xor in_data(68) xor in_data(70) xor in_data(72) xor in_data(74) xor in_data(75) xor in_data(76) xor in_data(77) xor in_data(79) xor in_data(80) xor in_data(82) xor in_data(83) xor in_data(89) xor in_data(90) xor in_data(92) xor in_data(95) xor in_data(97) xor in_data(100) xor in_data(101) xor in_data(109) xor in_data(113) xor in_data(117) xor in_data(118) xor in_data(119) xor in_data(120) xor in_data(122) xor in_data(123) xor in_data(124) xor in_data(127) xor in_data(133) xor in_data(134) xor in_data(135) xor in_data(137) xor in_data(138) xor in_data(139) xor in_data(141) xor in_data(143) xor in_data(144) xor in_data(148) xor in_data(150) xor in_data(151) xor in_data(152) xor in_data(153) xor in_data(157) xor in_data(159) xor in_data(163) xor in_data(166) xor in_data(170) xor in_data(172) xor in_data(173) xor in_data(176) xor in_data(177) xor in_data(179) xor in_data(181) xor in_data(182) xor in_data(184) xor in_data(185) xor in_data(187) xor in_data(188) xor in_data(189) xor in_data(190) xor in_data(191) xor in_data(192) xor in_data(194) xor in_data(195) xor in_data(199) xor in_data(200) xor in_data(204) xor in_data(213) xor in_data(214) xor in_data(215) xor in_data(216) xor in_data(221) xor in_data(223) xor in_data(226) xor in_data(228) xor in_data(229) xor in_data(230) xor in_data(237) xor in_data(239) xor in_data(240) xor in_data(242) xor in_data(245) xor in_data(246) xor in_data(248) xor in_data(249) xor in_data(250) xor in_data(251) xor in_data(254) xor in_data(256) xor in_data(261) xor in_data(262) xor in_data(267) xor in_data(268) xor in_data(269) xor in_data(274) xor in_data(275) xor in_data(277) xor in_data(278) xor in_data(279) xor in_data(281) xor in_data(282) xor in_data(285) xor in_data(288) xor in_data(291) xor in_data(293) xor in_data(295) xor in_data(298) xor in_data(303) xor in_data(308) xor in_data(309) xor in_data(310) xor in_data(311) xor in_data(312) xor in_data(313) xor in_data(314) xor in_data(315) xor in_data(316) xor in_data(318) xor in_data(320) xor in_data(321) xor in_data(322) xor in_data(323) xor in_data(324) xor in_data(327) xor in_data(328) xor in_data(329) xor in_data(332) xor in_data(334) xor in_data(335) xor in_data(336) xor in_data(337) xor in_data(338) xor in_data(339) xor in_data(340) xor in_data(343) xor in_data(346) xor in_data(347) xor in_data(348) xor in_data(350) xor in_data(351) xor in_data(353) xor in_data(355) xor in_data(356) xor in_data(357) xor in_data(360) xor in_data(361) xor in_data(362) xor in_data(363) xor in_data(364) xor in_data(366) xor in_data(367) xor in_data(368) xor in_data(369) xor in_data(370) xor in_data(372) xor in_data(378) xor in_data(381) xor in_data(383) xor in_data(384) xor in_data(386) xor in_data(387) xor in_data(388) xor in_data(392) xor in_data(393) xor in_data(394) xor in_data(397) xor in_data(398) xor in_data(402) xor in_data(403) xor in_data(404) xor in_data(405) xor in_data(406) xor in_data(412) xor in_data(414) xor in_data(416) xor in_data(418) xor in_data(420) xor in_data(421) xor in_data(424) xor in_data(426) xor in_data(428) xor in_data(429) xor in_data(430) xor in_data(432) xor in_data(436) xor in_data(437) xor in_data(439) xor in_data(441) xor in_data(443) xor in_data(447) xor in_data(448) xor in_data(449) xor in_data(451) xor in_data(454) xor in_data(457) xor in_data(458) xor in_data(460) xor in_data(464) xor in_data(466) xor in_data(468) xor in_data(469) xor in_data(471) xor in_data(473) xor in_data(476) xor in_data(477) xor in_data(478) xor in_data(479) xor in_data(480) xor in_data(481) xor in_data(485) xor in_data(486) xor in_data(488) xor in_data(489) xor in_data(491) xor in_data(496) xor in_data(498) xor in_data(499) xor in_data(500) xor in_data(502) xor in_data(503) xor in_data(504) xor in_data(505) xor in_data(507) xor in_data(509);

out_data(44)<= in_data(7) xor in_data(11) xor in_data(15) xor in_data(16) xor in_data(17) xor in_data(18) xor in_data(20) xor in_data(21) xor in_data(22) xor in_data(25) xor in_data(31) xor in_data(32) xor in_data(33) xor in_data(35) xor in_data(36) xor in_data(37) xor in_data(39) xor in_data(41) xor in_data(42) xor in_data(46) xor in_data(48) xor in_data(49) xor in_data(50) xor in_data(51) xor in_data(55) xor in_data(57) xor in_data(61) xor in_data(64) xor in_data(68) xor in_data(70) xor in_data(71) xor in_data(74) xor in_data(75) xor in_data(77) xor in_data(79) xor in_data(80) xor in_data(82) xor in_data(83) xor in_data(85) xor in_data(86) xor in_data(87) xor in_data(88) xor in_data(89) xor in_data(90) xor in_data(92) xor in_data(93) xor in_data(97) xor in_data(98) xor in_data(102) xor in_data(111) xor in_data(112) xor in_data(113) xor in_data(114) xor in_data(119) xor in_data(121) xor in_data(124) xor in_data(126) xor in_data(127) xor in_data(128) xor in_data(135) xor in_data(137) xor in_data(138) xor in_data(140) xor in_data(143) xor in_data(144) xor in_data(146) xor in_data(147) xor in_data(148) xor in_data(149) xor in_data(152) xor in_data(154) xor in_data(159) xor in_data(160) xor in_data(165) xor in_data(166) xor in_data(167) xor in_data(172) xor in_data(173) xor in_data(175) xor in_data(176) xor in_data(177) xor in_data(179) xor in_data(180) xor in_data(183) xor in_data(186) xor in_data(189) xor in_data(191) xor in_data(193) xor in_data(196) xor in_data(201) xor in_data(206) xor in_data(207) xor in_data(208) xor in_data(209) xor in_data(210) xor in_data(211) xor in_data(212) xor in_data(213) xor in_data(214) xor in_data(216) xor in_data(218) xor in_data(219) xor in_data(220) xor in_data(221) xor in_data(222) xor in_data(225) xor in_data(226) xor in_data(227) xor in_data(230) xor in_data(232) xor in_data(233) xor in_data(234) xor in_data(235) xor in_data(236) xor in_data(237) xor in_data(238) xor in_data(241) xor in_data(244) xor in_data(245) xor in_data(246) xor in_data(248) xor in_data(249) xor in_data(251) xor in_data(253) xor in_data(254) xor in_data(255) xor in_data(258) xor in_data(259) xor in_data(260) xor in_data(261) xor in_data(262) xor in_data(264) xor in_data(265) xor in_data(266) xor in_data(267) xor in_data(268) xor in_data(270) xor in_data(276) xor in_data(279) xor in_data(281) xor in_data(282) xor in_data(284) xor in_data(285) xor in_data(286) xor in_data(290) xor in_data(291) xor in_data(292) xor in_data(295) xor in_data(296) xor in_data(300) xor in_data(301) xor in_data(302) xor in_data(303) xor in_data(304) xor in_data(310) xor in_data(312) xor in_data(314) xor in_data(316) xor in_data(318) xor in_data(319) xor in_data(322) xor in_data(324) xor in_data(326) xor in_data(327) xor in_data(328) xor in_data(330) xor in_data(334) xor in_data(335) xor in_data(337) xor in_data(339) xor in_data(341) xor in_data(345) xor in_data(346) xor in_data(347) xor in_data(349) xor in_data(352) xor in_data(355) xor in_data(356) xor in_data(358) xor in_data(362) xor in_data(364) xor in_data(366) xor in_data(367) xor in_data(369) xor in_data(371) xor in_data(374) xor in_data(375) xor in_data(376) xor in_data(377) xor in_data(378) xor in_data(379) xor in_data(383) xor in_data(384) xor in_data(386) xor in_data(387) xor in_data(389) xor in_data(394) xor in_data(396) xor in_data(397) xor in_data(398) xor in_data(400) xor in_data(401) xor in_data(402) xor in_data(403) xor in_data(405) xor in_data(407) xor in_data(414) xor in_data(415) xor in_data(418) xor in_data(419) xor in_data(422) xor in_data(426) xor in_data(427) xor in_data(430) xor in_data(432) xor in_data(433) xor in_data(438) xor in_data(441) xor in_data(442) xor in_data(445) xor in_data(446) xor in_data(447) xor in_data(448) xor in_data(450) xor in_data(453) xor in_data(454) xor in_data(455) xor in_data(459) xor in_data(462) xor in_data(463) xor in_data(464) xor in_data(465) xor in_data(468) xor in_data(469) xor in_data(471) xor in_data(472) xor in_data(475) xor in_data(476) xor in_data(477) xor in_data(479) xor in_data(481) xor in_data(483) xor in_data(484) xor in_data(485) xor in_data(486) xor in_data(488) xor in_data(489) xor in_data(491) xor in_data(492) xor in_data(498) xor in_data(499) xor in_data(501) xor in_data(504) xor in_data(506) xor in_data(509) xor in_data(510);

out_data(45)<='0';

out_data(46)<='0';

out_data(47)<='0';

out_data(48)<='0';

out_data(49)<='0';

out_data(50)<='0';

out_data(51)<='0';

out_data(52)<='0';

out_data(53)<='0';

end;