library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.ALL;
package word_expander_package_for_D64_N113 is

    constant INPUT_WIDTH : integer := 64;
    constant OUTPUT_WIDTH : integer := 113;
    constant INPUT_ROM_ROWS : integer := 16;


    type ROM_type_expanded is array (0 to (INPUT_WIDTH*INPUT_ROM_ROWS-1)) of std_logic_vector((OUTPUT_WIDTH-1) downto 0);
    constant ROM_expanded : ROM_type_expanded := (
            "00000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000",
            "00000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "00001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111",
            "11111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "11111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000",
            "00000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "00000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111",
            "11111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "11111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111",
            "10000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "00000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000",
            "00000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "11111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111",
            "11111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "00000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000",
            "00000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "11111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111",
            "11111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "11000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000",
            "00000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "00000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111",
            "11111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "11111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000",
            "00000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "00000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001",
            "11111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "11111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111",
            "11100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "00000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000",
            "00000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "11111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
            "11111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "00000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000",
            "00000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111",
            "11111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "11110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000",
            "00000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "00000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111",
            "11111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "11111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000",
            "00000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "00000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000",
            "01111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "11111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111",
            "11111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "00000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000",
            "00000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "11111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
            "11111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "00000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000",
            "00000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "00111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111",
            "11111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "11111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000",
            "00000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "00000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111",
            "11111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "11111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110",
            "00000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "00000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000",
            "00011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "11111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111",
            "11111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "00000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000",
            "00000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "11111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111",
            "11111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000",
            "00000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "00001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111",
            "11111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "11111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000",
            "00000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "00000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111",
            "11111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "11111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111",
            "10000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "00000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000",
            "00000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "11111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111",
            "11111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "00000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000",
            "00000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "11111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111",
            "11111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "11000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000",
            "00000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "00000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111",
            "11111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "11111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000",
            "00000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "00000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001",
            "11111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "11111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111",
            "11100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "00000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000",
            "00000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "11111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
            "11111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "00000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000",
            "00000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111",
            "11111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "11110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000",
            "00000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "00000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111",
            "11111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "11111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000",
            "00000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "00000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000",
            "01111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "11111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111",
            "11111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "00000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000",
            "00000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "11111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
            "11111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "00000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000",
            "00000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "00111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111",
            "11111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "11111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000",
            "00000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "00000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111",
            "11111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "11111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110",
            "00000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "00000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000",
            "00011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "11111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111",
            "11111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "00000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000",
            "00000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "11111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111",
            "11111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000",
            "00000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "00001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111",
            "11111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "11111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000",
            "00000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "00000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111",
            "11111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "11111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111",
            "10000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "00000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000",
            "00000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "11111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111",
            "11111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "00000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000",
            "00000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "11111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111",
            "11111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "11000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000",
            "00000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "00000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111",
            "11111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "11111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000",
            "00000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "00000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001",
            "11111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "11111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111",
            "11100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "00000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000",
            "00000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "11111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
            "11111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "00000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000",
            "00000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111",
            "11111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "11110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000",
            "00000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "00000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111",
            "11111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "11111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000",
            "00000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "00000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000",
            "01111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "11111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111",
            "11111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "00000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000",
            "00000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "11111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
            "11111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "00000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000",
            "00000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "00111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111",
            "11111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "11111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000",
            "00000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "00000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111",
            "11111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "11111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110",
            "00000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "00000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000",
            "00011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "11111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111",
            "11111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "00000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000",
            "00000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "11111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111",
            "11111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000",
            "00000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "00001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111",
            "11111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "11111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000",
            "00000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "00000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111",
            "11111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "11111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111",
            "10000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "00000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000",
            "00000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "11111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111",
            "11111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "00000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000",
            "00000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "11111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111",
            "11111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "11000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000",
            "00000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "00000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111",
            "11111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "11111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000",
            "00000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "00000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001",
            "11111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "11111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111",
            "11100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "00000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000",
            "00000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "11111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
            "11111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "00000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000",
            "00000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111",
            "11111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "11110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000",
            "00000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "00000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111",
            "11111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "11111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000",
            "00000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "00000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000",
            "01111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "11111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111",
            "11111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "00000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000",
            "00000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "11111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
            "11111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "00000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000",
            "00000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "00111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111",
            "11111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "11111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000",
            "00000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "00000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111",
            "11111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "11111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110",
            "00000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "00000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000",
            "00011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "11111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111",
            "11111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "00000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000",
            "00000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "11111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111",
            "11111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000",
            "00000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "00001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111",
            "11111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "11111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000",
            "00000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "00000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111",
            "11111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "11111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111",
            "10000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "00000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000",
            "00000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "11111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111",
            "11111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "00000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000",
            "00000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "11111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111",
            "11111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "11000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000",
            "00000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "00000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111",
            "11111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "11111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000",
            "00000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "00000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001",
            "11111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "11111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111",
            "11100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "00000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000",
            "00000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "11111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
            "11111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "00000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000",
            "00000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111",
            "11111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "11110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000",
            "00000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "00000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111",
            "11111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "11111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000",
            "00000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "00000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000",
            "01111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "11111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111",
            "11111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "00000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000",
            "00000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "11111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
            "11111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "00000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000",
            "00000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "00111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111",
            "11111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "11111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000",
            "00000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "00000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111",
            "11111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "11111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110",
            "00000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "00000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000",
            "00011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "11111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111",
            "11111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "00000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000",
            "00000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "11111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111",
            "11111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000",
            "00000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "00001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111",
            "11111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "11111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000",
            "00000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "00000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111",
            "11111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "11111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111",
            "10000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "00000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000",
            "00000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "11111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111",
            "11111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "00000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000",
            "00000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "11111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111",
            "11111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "11000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000",
            "00000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "00000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111",
            "11111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "11111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000",
            "00000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "00000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001",
            "11111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "11111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111",
            "11100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "00000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000",
            "00000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "11111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
            "11111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "00000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000",
            "00000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111",
            "11111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "11110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000",
            "00000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "00000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111",
            "11111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "11111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000",
            "00000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "00000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000",
            "01111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "11111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111",
            "11111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "00000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000",
            "00000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "11111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
            "11111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "00000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000",
            "00000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "00111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111",
            "11111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "11111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000",
            "00000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "00000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111",
            "11111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "11111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110",
            "00000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "00000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000",
            "00011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "11111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111",
            "11111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "00000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000",
            "00000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "11111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111",
            "11111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000",
            "00000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "00001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111",
            "11111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "11111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000",
            "00000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "00000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111",
            "11111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "11111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111",
            "10000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "00000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000",
            "00000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "11111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111",
            "11111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "00000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000",
            "00000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "11111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111",
            "11111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "11000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000",
            "00000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "00000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111",
            "11111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "11111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000",
            "00000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "00000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001",
            "11111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "11111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111",
            "11100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "00000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000",
            "00000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "11111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
            "11111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "00000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000",
            "00000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111",
            "11111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "11110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000",
            "00000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "00000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111",
            "11111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "11111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000",
            "00000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "00000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000",
            "01111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "11111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111",
            "11111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "00000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000",
            "00000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "11111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
            "11111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "00000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000",
            "00000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "00111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111",
            "11111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "11111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000",
            "00000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "00000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111",
            "11111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "11111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110",
            "00000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "00000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000",
            "00011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "11111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111",
            "11111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "00000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000",
            "00000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "11111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111",
            "11111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000",
            "00000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000",
            "00001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111",
            "11111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
            "11111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000",
            "00000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000",
            "00000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111",
            "11111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111",
            "11111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111",
            "10000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000",
            "00000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000",
            "00000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111",
            "11111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111",
            "11111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000",
            "00000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000",
            "00000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011",
            "11111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111",
            "11111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111",
            "11000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000",
            "00000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000",
            "00000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111",
            "11111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
            "11111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000",
            "00000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000",
            "00000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001",
            "11111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111",
            "11111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111",
            "11100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000",
            "00000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000",
            "00000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
            "11111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
            "11111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000",
            "00000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000",
            "00000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111",
            "11111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
            "11110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000",
            "00000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000",
            "00000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111",
            "11111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
            "11111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000",
            "00000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000",
            "00000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000",
            "01111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111",
            "11111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111",
            "11111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000",
            "00000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000",
            "00000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111",
            "11111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
            "11111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100",
            "00000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000",
            "00000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000",
            "00111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111",
            "11111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
            "11111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000",
            "00000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000",
            "00000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111",
            "11111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
            "11111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110",
            "00000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000",
            "00000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000",
            "00011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111",
            "11111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111",
            "11111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
            "00000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000",
            "00000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000",
            "00000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000",
            "11111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111",
            "11111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111",
            "11111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
            "00000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111"
    );

    type ROM_type_data is array (0 to (INPUT_ROM_ROWS-1)) of std_logic_vector((INPUT_WIDTH-1) downto 0);
    constant ROM_data : ROM_type_data := (
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000"
    );

    function ROM_send_data(index : integer) return std_logic_vector;    function ROM_D64_N113(index : integer) return std_logic_vector;

end word_expander_package_for_D64_N113;

package body word_expander_package_for_D64_N113 is

    function ROM_send_data(index : integer) return std_logic_vector is
    begin
        return ROM_data(index);
    end ROM_send_data;


    function ROM_D64_N113(index : integer) return std_logic_vector is
    begin
        return ROM_expanded(index);
    end ROM_D64_N113;


end word_expander_package_for_D64_N113;