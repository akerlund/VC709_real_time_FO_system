library ieee;
use ieee.std_logic_1164.all;
entity chien is
    port(
        a_1     :    in  std_logic_vector(9 downto 0);
        a_2     :    in  std_logic_vector(9 downto 0);
        a_3     :    in  std_logic_vector(9 downto 0);
        a_4     :    in  std_logic_vector(9 downto 0);
        E     :    out std_logic_vector(1022 downto 0)
);
end entity;

architecture arch of chien is
    signal mulr_1_1 : std_logic_vector(9 downto 0);
    signal mulr_2_1 : std_logic_vector(9 downto 0);
    signal mulr_3_1 : std_logic_vector(9 downto 0);
    signal mulr_4_1 : std_logic_vector(9 downto 0);
    signal mulr_1_2 : std_logic_vector(9 downto 0);
    signal mulr_2_2 : std_logic_vector(9 downto 0);
    signal mulr_3_2 : std_logic_vector(9 downto 0);
    signal mulr_4_2 : std_logic_vector(9 downto 0);
    signal mulr_1_3 : std_logic_vector(9 downto 0);
    signal mulr_2_3 : std_logic_vector(9 downto 0);
    signal mulr_3_3 : std_logic_vector(9 downto 0);
    signal mulr_4_3 : std_logic_vector(9 downto 0);
    signal mulr_1_4 : std_logic_vector(9 downto 0);
    signal mulr_2_4 : std_logic_vector(9 downto 0);
    signal mulr_3_4 : std_logic_vector(9 downto 0);
    signal mulr_4_4 : std_logic_vector(9 downto 0);
    signal mulr_1_5 : std_logic_vector(9 downto 0);
    signal mulr_2_5 : std_logic_vector(9 downto 0);
    signal mulr_3_5 : std_logic_vector(9 downto 0);
    signal mulr_4_5 : std_logic_vector(9 downto 0);
    signal mulr_1_6 : std_logic_vector(9 downto 0);
    signal mulr_2_6 : std_logic_vector(9 downto 0);
    signal mulr_3_6 : std_logic_vector(9 downto 0);
    signal mulr_4_6 : std_logic_vector(9 downto 0);
    signal mulr_1_7 : std_logic_vector(9 downto 0);
    signal mulr_2_7 : std_logic_vector(9 downto 0);
    signal mulr_3_7 : std_logic_vector(9 downto 0);
    signal mulr_4_7 : std_logic_vector(9 downto 0);
    signal mulr_1_8 : std_logic_vector(9 downto 0);
    signal mulr_2_8 : std_logic_vector(9 downto 0);
    signal mulr_3_8 : std_logic_vector(9 downto 0);
    signal mulr_4_8 : std_logic_vector(9 downto 0);
    signal mulr_1_9 : std_logic_vector(9 downto 0);
    signal mulr_2_9 : std_logic_vector(9 downto 0);
    signal mulr_3_9 : std_logic_vector(9 downto 0);
    signal mulr_4_9 : std_logic_vector(9 downto 0);
    signal mulr_1_10 : std_logic_vector(9 downto 0);
    signal mulr_2_10 : std_logic_vector(9 downto 0);
    signal mulr_3_10 : std_logic_vector(9 downto 0);
    signal mulr_4_10 : std_logic_vector(9 downto 0);
    signal mulr_1_11 : std_logic_vector(9 downto 0);
    signal mulr_2_11 : std_logic_vector(9 downto 0);
    signal mulr_3_11 : std_logic_vector(9 downto 0);
    signal mulr_4_11 : std_logic_vector(9 downto 0);
    signal mulr_1_12 : std_logic_vector(9 downto 0);
    signal mulr_2_12 : std_logic_vector(9 downto 0);
    signal mulr_3_12 : std_logic_vector(9 downto 0);
    signal mulr_4_12 : std_logic_vector(9 downto 0);
    signal mulr_1_13 : std_logic_vector(9 downto 0);
    signal mulr_2_13 : std_logic_vector(9 downto 0);
    signal mulr_3_13 : std_logic_vector(9 downto 0);
    signal mulr_4_13 : std_logic_vector(9 downto 0);
    signal mulr_1_14 : std_logic_vector(9 downto 0);
    signal mulr_2_14 : std_logic_vector(9 downto 0);
    signal mulr_3_14 : std_logic_vector(9 downto 0);
    signal mulr_4_14 : std_logic_vector(9 downto 0);
    signal mulr_1_15 : std_logic_vector(9 downto 0);
    signal mulr_2_15 : std_logic_vector(9 downto 0);
    signal mulr_3_15 : std_logic_vector(9 downto 0);
    signal mulr_4_15 : std_logic_vector(9 downto 0);
    signal mulr_1_16 : std_logic_vector(9 downto 0);
    signal mulr_2_16 : std_logic_vector(9 downto 0);
    signal mulr_3_16 : std_logic_vector(9 downto 0);
    signal mulr_4_16 : std_logic_vector(9 downto 0);
    signal mulr_1_17 : std_logic_vector(9 downto 0);
    signal mulr_2_17 : std_logic_vector(9 downto 0);
    signal mulr_3_17 : std_logic_vector(9 downto 0);
    signal mulr_4_17 : std_logic_vector(9 downto 0);
    signal mulr_1_18 : std_logic_vector(9 downto 0);
    signal mulr_2_18 : std_logic_vector(9 downto 0);
    signal mulr_3_18 : std_logic_vector(9 downto 0);
    signal mulr_4_18 : std_logic_vector(9 downto 0);
    signal mulr_1_19 : std_logic_vector(9 downto 0);
    signal mulr_2_19 : std_logic_vector(9 downto 0);
    signal mulr_3_19 : std_logic_vector(9 downto 0);
    signal mulr_4_19 : std_logic_vector(9 downto 0);
    signal mulr_1_20 : std_logic_vector(9 downto 0);
    signal mulr_2_20 : std_logic_vector(9 downto 0);
    signal mulr_3_20 : std_logic_vector(9 downto 0);
    signal mulr_4_20 : std_logic_vector(9 downto 0);
    signal mulr_1_21 : std_logic_vector(9 downto 0);
    signal mulr_2_21 : std_logic_vector(9 downto 0);
    signal mulr_3_21 : std_logic_vector(9 downto 0);
    signal mulr_4_21 : std_logic_vector(9 downto 0);
    signal mulr_1_22 : std_logic_vector(9 downto 0);
    signal mulr_2_22 : std_logic_vector(9 downto 0);
    signal mulr_3_22 : std_logic_vector(9 downto 0);
    signal mulr_4_22 : std_logic_vector(9 downto 0);
    signal mulr_1_23 : std_logic_vector(9 downto 0);
    signal mulr_2_23 : std_logic_vector(9 downto 0);
    signal mulr_3_23 : std_logic_vector(9 downto 0);
    signal mulr_4_23 : std_logic_vector(9 downto 0);
    signal mulr_1_24 : std_logic_vector(9 downto 0);
    signal mulr_2_24 : std_logic_vector(9 downto 0);
    signal mulr_3_24 : std_logic_vector(9 downto 0);
    signal mulr_4_24 : std_logic_vector(9 downto 0);
    signal mulr_1_25 : std_logic_vector(9 downto 0);
    signal mulr_2_25 : std_logic_vector(9 downto 0);
    signal mulr_3_25 : std_logic_vector(9 downto 0);
    signal mulr_4_25 : std_logic_vector(9 downto 0);
    signal mulr_1_26 : std_logic_vector(9 downto 0);
    signal mulr_2_26 : std_logic_vector(9 downto 0);
    signal mulr_3_26 : std_logic_vector(9 downto 0);
    signal mulr_4_26 : std_logic_vector(9 downto 0);
    signal mulr_1_27 : std_logic_vector(9 downto 0);
    signal mulr_2_27 : std_logic_vector(9 downto 0);
    signal mulr_3_27 : std_logic_vector(9 downto 0);
    signal mulr_4_27 : std_logic_vector(9 downto 0);
    signal mulr_1_28 : std_logic_vector(9 downto 0);
    signal mulr_2_28 : std_logic_vector(9 downto 0);
    signal mulr_3_28 : std_logic_vector(9 downto 0);
    signal mulr_4_28 : std_logic_vector(9 downto 0);
    signal mulr_1_29 : std_logic_vector(9 downto 0);
    signal mulr_2_29 : std_logic_vector(9 downto 0);
    signal mulr_3_29 : std_logic_vector(9 downto 0);
    signal mulr_4_29 : std_logic_vector(9 downto 0);
    signal mulr_1_30 : std_logic_vector(9 downto 0);
    signal mulr_2_30 : std_logic_vector(9 downto 0);
    signal mulr_3_30 : std_logic_vector(9 downto 0);
    signal mulr_4_30 : std_logic_vector(9 downto 0);
    signal mulr_1_31 : std_logic_vector(9 downto 0);
    signal mulr_2_31 : std_logic_vector(9 downto 0);
    signal mulr_3_31 : std_logic_vector(9 downto 0);
    signal mulr_4_31 : std_logic_vector(9 downto 0);
    signal mulr_1_32 : std_logic_vector(9 downto 0);
    signal mulr_2_32 : std_logic_vector(9 downto 0);
    signal mulr_3_32 : std_logic_vector(9 downto 0);
    signal mulr_4_32 : std_logic_vector(9 downto 0);
    signal mulr_1_33 : std_logic_vector(9 downto 0);
    signal mulr_2_33 : std_logic_vector(9 downto 0);
    signal mulr_3_33 : std_logic_vector(9 downto 0);
    signal mulr_4_33 : std_logic_vector(9 downto 0);
    signal mulr_1_34 : std_logic_vector(9 downto 0);
    signal mulr_2_34 : std_logic_vector(9 downto 0);
    signal mulr_3_34 : std_logic_vector(9 downto 0);
    signal mulr_4_34 : std_logic_vector(9 downto 0);
    signal mulr_1_35 : std_logic_vector(9 downto 0);
    signal mulr_2_35 : std_logic_vector(9 downto 0);
    signal mulr_3_35 : std_logic_vector(9 downto 0);
    signal mulr_4_35 : std_logic_vector(9 downto 0);
    signal mulr_1_36 : std_logic_vector(9 downto 0);
    signal mulr_2_36 : std_logic_vector(9 downto 0);
    signal mulr_3_36 : std_logic_vector(9 downto 0);
    signal mulr_4_36 : std_logic_vector(9 downto 0);
    signal mulr_1_37 : std_logic_vector(9 downto 0);
    signal mulr_2_37 : std_logic_vector(9 downto 0);
    signal mulr_3_37 : std_logic_vector(9 downto 0);
    signal mulr_4_37 : std_logic_vector(9 downto 0);
    signal mulr_1_38 : std_logic_vector(9 downto 0);
    signal mulr_2_38 : std_logic_vector(9 downto 0);
    signal mulr_3_38 : std_logic_vector(9 downto 0);
    signal mulr_4_38 : std_logic_vector(9 downto 0);
    signal mulr_1_39 : std_logic_vector(9 downto 0);
    signal mulr_2_39 : std_logic_vector(9 downto 0);
    signal mulr_3_39 : std_logic_vector(9 downto 0);
    signal mulr_4_39 : std_logic_vector(9 downto 0);
    signal mulr_1_40 : std_logic_vector(9 downto 0);
    signal mulr_2_40 : std_logic_vector(9 downto 0);
    signal mulr_3_40 : std_logic_vector(9 downto 0);
    signal mulr_4_40 : std_logic_vector(9 downto 0);
    signal mulr_1_41 : std_logic_vector(9 downto 0);
    signal mulr_2_41 : std_logic_vector(9 downto 0);
    signal mulr_3_41 : std_logic_vector(9 downto 0);
    signal mulr_4_41 : std_logic_vector(9 downto 0);
    signal mulr_1_42 : std_logic_vector(9 downto 0);
    signal mulr_2_42 : std_logic_vector(9 downto 0);
    signal mulr_3_42 : std_logic_vector(9 downto 0);
    signal mulr_4_42 : std_logic_vector(9 downto 0);
    signal mulr_1_43 : std_logic_vector(9 downto 0);
    signal mulr_2_43 : std_logic_vector(9 downto 0);
    signal mulr_3_43 : std_logic_vector(9 downto 0);
    signal mulr_4_43 : std_logic_vector(9 downto 0);
    signal mulr_1_44 : std_logic_vector(9 downto 0);
    signal mulr_2_44 : std_logic_vector(9 downto 0);
    signal mulr_3_44 : std_logic_vector(9 downto 0);
    signal mulr_4_44 : std_logic_vector(9 downto 0);
    signal mulr_1_45 : std_logic_vector(9 downto 0);
    signal mulr_2_45 : std_logic_vector(9 downto 0);
    signal mulr_3_45 : std_logic_vector(9 downto 0);
    signal mulr_4_45 : std_logic_vector(9 downto 0);
    signal mulr_1_46 : std_logic_vector(9 downto 0);
    signal mulr_2_46 : std_logic_vector(9 downto 0);
    signal mulr_3_46 : std_logic_vector(9 downto 0);
    signal mulr_4_46 : std_logic_vector(9 downto 0);
    signal mulr_1_47 : std_logic_vector(9 downto 0);
    signal mulr_2_47 : std_logic_vector(9 downto 0);
    signal mulr_3_47 : std_logic_vector(9 downto 0);
    signal mulr_4_47 : std_logic_vector(9 downto 0);
    signal mulr_1_48 : std_logic_vector(9 downto 0);
    signal mulr_2_48 : std_logic_vector(9 downto 0);
    signal mulr_3_48 : std_logic_vector(9 downto 0);
    signal mulr_4_48 : std_logic_vector(9 downto 0);
    signal mulr_1_49 : std_logic_vector(9 downto 0);
    signal mulr_2_49 : std_logic_vector(9 downto 0);
    signal mulr_3_49 : std_logic_vector(9 downto 0);
    signal mulr_4_49 : std_logic_vector(9 downto 0);
    signal mulr_1_50 : std_logic_vector(9 downto 0);
    signal mulr_2_50 : std_logic_vector(9 downto 0);
    signal mulr_3_50 : std_logic_vector(9 downto 0);
    signal mulr_4_50 : std_logic_vector(9 downto 0);
    signal mulr_1_51 : std_logic_vector(9 downto 0);
    signal mulr_2_51 : std_logic_vector(9 downto 0);
    signal mulr_3_51 : std_logic_vector(9 downto 0);
    signal mulr_4_51 : std_logic_vector(9 downto 0);
    signal mulr_1_52 : std_logic_vector(9 downto 0);
    signal mulr_2_52 : std_logic_vector(9 downto 0);
    signal mulr_3_52 : std_logic_vector(9 downto 0);
    signal mulr_4_52 : std_logic_vector(9 downto 0);
    signal mulr_1_53 : std_logic_vector(9 downto 0);
    signal mulr_2_53 : std_logic_vector(9 downto 0);
    signal mulr_3_53 : std_logic_vector(9 downto 0);
    signal mulr_4_53 : std_logic_vector(9 downto 0);
    signal mulr_1_54 : std_logic_vector(9 downto 0);
    signal mulr_2_54 : std_logic_vector(9 downto 0);
    signal mulr_3_54 : std_logic_vector(9 downto 0);
    signal mulr_4_54 : std_logic_vector(9 downto 0);
    signal mulr_1_55 : std_logic_vector(9 downto 0);
    signal mulr_2_55 : std_logic_vector(9 downto 0);
    signal mulr_3_55 : std_logic_vector(9 downto 0);
    signal mulr_4_55 : std_logic_vector(9 downto 0);
    signal mulr_1_56 : std_logic_vector(9 downto 0);
    signal mulr_2_56 : std_logic_vector(9 downto 0);
    signal mulr_3_56 : std_logic_vector(9 downto 0);
    signal mulr_4_56 : std_logic_vector(9 downto 0);
    signal mulr_1_57 : std_logic_vector(9 downto 0);
    signal mulr_2_57 : std_logic_vector(9 downto 0);
    signal mulr_3_57 : std_logic_vector(9 downto 0);
    signal mulr_4_57 : std_logic_vector(9 downto 0);
    signal mulr_1_58 : std_logic_vector(9 downto 0);
    signal mulr_2_58 : std_logic_vector(9 downto 0);
    signal mulr_3_58 : std_logic_vector(9 downto 0);
    signal mulr_4_58 : std_logic_vector(9 downto 0);
    signal mulr_1_59 : std_logic_vector(9 downto 0);
    signal mulr_2_59 : std_logic_vector(9 downto 0);
    signal mulr_3_59 : std_logic_vector(9 downto 0);
    signal mulr_4_59 : std_logic_vector(9 downto 0);
    signal mulr_1_60 : std_logic_vector(9 downto 0);
    signal mulr_2_60 : std_logic_vector(9 downto 0);
    signal mulr_3_60 : std_logic_vector(9 downto 0);
    signal mulr_4_60 : std_logic_vector(9 downto 0);
    signal mulr_1_61 : std_logic_vector(9 downto 0);
    signal mulr_2_61 : std_logic_vector(9 downto 0);
    signal mulr_3_61 : std_logic_vector(9 downto 0);
    signal mulr_4_61 : std_logic_vector(9 downto 0);
    signal mulr_1_62 : std_logic_vector(9 downto 0);
    signal mulr_2_62 : std_logic_vector(9 downto 0);
    signal mulr_3_62 : std_logic_vector(9 downto 0);
    signal mulr_4_62 : std_logic_vector(9 downto 0);
    signal mulr_1_63 : std_logic_vector(9 downto 0);
    signal mulr_2_63 : std_logic_vector(9 downto 0);
    signal mulr_3_63 : std_logic_vector(9 downto 0);
    signal mulr_4_63 : std_logic_vector(9 downto 0);
    signal mulr_1_64 : std_logic_vector(9 downto 0);
    signal mulr_2_64 : std_logic_vector(9 downto 0);
    signal mulr_3_64 : std_logic_vector(9 downto 0);
    signal mulr_4_64 : std_logic_vector(9 downto 0);
    signal mulr_1_65 : std_logic_vector(9 downto 0);
    signal mulr_2_65 : std_logic_vector(9 downto 0);
    signal mulr_3_65 : std_logic_vector(9 downto 0);
    signal mulr_4_65 : std_logic_vector(9 downto 0);
    signal mulr_1_66 : std_logic_vector(9 downto 0);
    signal mulr_2_66 : std_logic_vector(9 downto 0);
    signal mulr_3_66 : std_logic_vector(9 downto 0);
    signal mulr_4_66 : std_logic_vector(9 downto 0);
    signal mulr_1_67 : std_logic_vector(9 downto 0);
    signal mulr_2_67 : std_logic_vector(9 downto 0);
    signal mulr_3_67 : std_logic_vector(9 downto 0);
    signal mulr_4_67 : std_logic_vector(9 downto 0);
    signal mulr_1_68 : std_logic_vector(9 downto 0);
    signal mulr_2_68 : std_logic_vector(9 downto 0);
    signal mulr_3_68 : std_logic_vector(9 downto 0);
    signal mulr_4_68 : std_logic_vector(9 downto 0);
    signal mulr_1_69 : std_logic_vector(9 downto 0);
    signal mulr_2_69 : std_logic_vector(9 downto 0);
    signal mulr_3_69 : std_logic_vector(9 downto 0);
    signal mulr_4_69 : std_logic_vector(9 downto 0);
    signal mulr_1_70 : std_logic_vector(9 downto 0);
    signal mulr_2_70 : std_logic_vector(9 downto 0);
    signal mulr_3_70 : std_logic_vector(9 downto 0);
    signal mulr_4_70 : std_logic_vector(9 downto 0);
    signal mulr_1_71 : std_logic_vector(9 downto 0);
    signal mulr_2_71 : std_logic_vector(9 downto 0);
    signal mulr_3_71 : std_logic_vector(9 downto 0);
    signal mulr_4_71 : std_logic_vector(9 downto 0);
    signal mulr_1_72 : std_logic_vector(9 downto 0);
    signal mulr_2_72 : std_logic_vector(9 downto 0);
    signal mulr_3_72 : std_logic_vector(9 downto 0);
    signal mulr_4_72 : std_logic_vector(9 downto 0);
    signal mulr_1_73 : std_logic_vector(9 downto 0);
    signal mulr_2_73 : std_logic_vector(9 downto 0);
    signal mulr_3_73 : std_logic_vector(9 downto 0);
    signal mulr_4_73 : std_logic_vector(9 downto 0);
    signal mulr_1_74 : std_logic_vector(9 downto 0);
    signal mulr_2_74 : std_logic_vector(9 downto 0);
    signal mulr_3_74 : std_logic_vector(9 downto 0);
    signal mulr_4_74 : std_logic_vector(9 downto 0);
    signal mulr_1_75 : std_logic_vector(9 downto 0);
    signal mulr_2_75 : std_logic_vector(9 downto 0);
    signal mulr_3_75 : std_logic_vector(9 downto 0);
    signal mulr_4_75 : std_logic_vector(9 downto 0);
    signal mulr_1_76 : std_logic_vector(9 downto 0);
    signal mulr_2_76 : std_logic_vector(9 downto 0);
    signal mulr_3_76 : std_logic_vector(9 downto 0);
    signal mulr_4_76 : std_logic_vector(9 downto 0);
    signal mulr_1_77 : std_logic_vector(9 downto 0);
    signal mulr_2_77 : std_logic_vector(9 downto 0);
    signal mulr_3_77 : std_logic_vector(9 downto 0);
    signal mulr_4_77 : std_logic_vector(9 downto 0);
    signal mulr_1_78 : std_logic_vector(9 downto 0);
    signal mulr_2_78 : std_logic_vector(9 downto 0);
    signal mulr_3_78 : std_logic_vector(9 downto 0);
    signal mulr_4_78 : std_logic_vector(9 downto 0);
    signal mulr_1_79 : std_logic_vector(9 downto 0);
    signal mulr_2_79 : std_logic_vector(9 downto 0);
    signal mulr_3_79 : std_logic_vector(9 downto 0);
    signal mulr_4_79 : std_logic_vector(9 downto 0);
    signal mulr_1_80 : std_logic_vector(9 downto 0);
    signal mulr_2_80 : std_logic_vector(9 downto 0);
    signal mulr_3_80 : std_logic_vector(9 downto 0);
    signal mulr_4_80 : std_logic_vector(9 downto 0);
    signal mulr_1_81 : std_logic_vector(9 downto 0);
    signal mulr_2_81 : std_logic_vector(9 downto 0);
    signal mulr_3_81 : std_logic_vector(9 downto 0);
    signal mulr_4_81 : std_logic_vector(9 downto 0);
    signal mulr_1_82 : std_logic_vector(9 downto 0);
    signal mulr_2_82 : std_logic_vector(9 downto 0);
    signal mulr_3_82 : std_logic_vector(9 downto 0);
    signal mulr_4_82 : std_logic_vector(9 downto 0);
    signal mulr_1_83 : std_logic_vector(9 downto 0);
    signal mulr_2_83 : std_logic_vector(9 downto 0);
    signal mulr_3_83 : std_logic_vector(9 downto 0);
    signal mulr_4_83 : std_logic_vector(9 downto 0);
    signal mulr_1_84 : std_logic_vector(9 downto 0);
    signal mulr_2_84 : std_logic_vector(9 downto 0);
    signal mulr_3_84 : std_logic_vector(9 downto 0);
    signal mulr_4_84 : std_logic_vector(9 downto 0);
    signal mulr_1_85 : std_logic_vector(9 downto 0);
    signal mulr_2_85 : std_logic_vector(9 downto 0);
    signal mulr_3_85 : std_logic_vector(9 downto 0);
    signal mulr_4_85 : std_logic_vector(9 downto 0);
    signal mulr_1_86 : std_logic_vector(9 downto 0);
    signal mulr_2_86 : std_logic_vector(9 downto 0);
    signal mulr_3_86 : std_logic_vector(9 downto 0);
    signal mulr_4_86 : std_logic_vector(9 downto 0);
    signal mulr_1_87 : std_logic_vector(9 downto 0);
    signal mulr_2_87 : std_logic_vector(9 downto 0);
    signal mulr_3_87 : std_logic_vector(9 downto 0);
    signal mulr_4_87 : std_logic_vector(9 downto 0);
    signal mulr_1_88 : std_logic_vector(9 downto 0);
    signal mulr_2_88 : std_logic_vector(9 downto 0);
    signal mulr_3_88 : std_logic_vector(9 downto 0);
    signal mulr_4_88 : std_logic_vector(9 downto 0);
    signal mulr_1_89 : std_logic_vector(9 downto 0);
    signal mulr_2_89 : std_logic_vector(9 downto 0);
    signal mulr_3_89 : std_logic_vector(9 downto 0);
    signal mulr_4_89 : std_logic_vector(9 downto 0);
    signal mulr_1_90 : std_logic_vector(9 downto 0);
    signal mulr_2_90 : std_logic_vector(9 downto 0);
    signal mulr_3_90 : std_logic_vector(9 downto 0);
    signal mulr_4_90 : std_logic_vector(9 downto 0);
    signal mulr_1_91 : std_logic_vector(9 downto 0);
    signal mulr_2_91 : std_logic_vector(9 downto 0);
    signal mulr_3_91 : std_logic_vector(9 downto 0);
    signal mulr_4_91 : std_logic_vector(9 downto 0);
    signal mulr_1_92 : std_logic_vector(9 downto 0);
    signal mulr_2_92 : std_logic_vector(9 downto 0);
    signal mulr_3_92 : std_logic_vector(9 downto 0);
    signal mulr_4_92 : std_logic_vector(9 downto 0);
    signal mulr_1_93 : std_logic_vector(9 downto 0);
    signal mulr_2_93 : std_logic_vector(9 downto 0);
    signal mulr_3_93 : std_logic_vector(9 downto 0);
    signal mulr_4_93 : std_logic_vector(9 downto 0);
    signal mulr_1_94 : std_logic_vector(9 downto 0);
    signal mulr_2_94 : std_logic_vector(9 downto 0);
    signal mulr_3_94 : std_logic_vector(9 downto 0);
    signal mulr_4_94 : std_logic_vector(9 downto 0);
    signal mulr_1_95 : std_logic_vector(9 downto 0);
    signal mulr_2_95 : std_logic_vector(9 downto 0);
    signal mulr_3_95 : std_logic_vector(9 downto 0);
    signal mulr_4_95 : std_logic_vector(9 downto 0);
    signal mulr_1_96 : std_logic_vector(9 downto 0);
    signal mulr_2_96 : std_logic_vector(9 downto 0);
    signal mulr_3_96 : std_logic_vector(9 downto 0);
    signal mulr_4_96 : std_logic_vector(9 downto 0);
    signal mulr_1_97 : std_logic_vector(9 downto 0);
    signal mulr_2_97 : std_logic_vector(9 downto 0);
    signal mulr_3_97 : std_logic_vector(9 downto 0);
    signal mulr_4_97 : std_logic_vector(9 downto 0);
    signal mulr_1_98 : std_logic_vector(9 downto 0);
    signal mulr_2_98 : std_logic_vector(9 downto 0);
    signal mulr_3_98 : std_logic_vector(9 downto 0);
    signal mulr_4_98 : std_logic_vector(9 downto 0);
    signal mulr_1_99 : std_logic_vector(9 downto 0);
    signal mulr_2_99 : std_logic_vector(9 downto 0);
    signal mulr_3_99 : std_logic_vector(9 downto 0);
    signal mulr_4_99 : std_logic_vector(9 downto 0);
    signal mulr_1_100 : std_logic_vector(9 downto 0);
    signal mulr_2_100 : std_logic_vector(9 downto 0);
    signal mulr_3_100 : std_logic_vector(9 downto 0);
    signal mulr_4_100 : std_logic_vector(9 downto 0);
    signal mulr_1_101 : std_logic_vector(9 downto 0);
    signal mulr_2_101 : std_logic_vector(9 downto 0);
    signal mulr_3_101 : std_logic_vector(9 downto 0);
    signal mulr_4_101 : std_logic_vector(9 downto 0);
    signal mulr_1_102 : std_logic_vector(9 downto 0);
    signal mulr_2_102 : std_logic_vector(9 downto 0);
    signal mulr_3_102 : std_logic_vector(9 downto 0);
    signal mulr_4_102 : std_logic_vector(9 downto 0);
    signal mulr_1_103 : std_logic_vector(9 downto 0);
    signal mulr_2_103 : std_logic_vector(9 downto 0);
    signal mulr_3_103 : std_logic_vector(9 downto 0);
    signal mulr_4_103 : std_logic_vector(9 downto 0);
    signal mulr_1_104 : std_logic_vector(9 downto 0);
    signal mulr_2_104 : std_logic_vector(9 downto 0);
    signal mulr_3_104 : std_logic_vector(9 downto 0);
    signal mulr_4_104 : std_logic_vector(9 downto 0);
    signal mulr_1_105 : std_logic_vector(9 downto 0);
    signal mulr_2_105 : std_logic_vector(9 downto 0);
    signal mulr_3_105 : std_logic_vector(9 downto 0);
    signal mulr_4_105 : std_logic_vector(9 downto 0);
    signal mulr_1_106 : std_logic_vector(9 downto 0);
    signal mulr_2_106 : std_logic_vector(9 downto 0);
    signal mulr_3_106 : std_logic_vector(9 downto 0);
    signal mulr_4_106 : std_logic_vector(9 downto 0);
    signal mulr_1_107 : std_logic_vector(9 downto 0);
    signal mulr_2_107 : std_logic_vector(9 downto 0);
    signal mulr_3_107 : std_logic_vector(9 downto 0);
    signal mulr_4_107 : std_logic_vector(9 downto 0);
    signal mulr_1_108 : std_logic_vector(9 downto 0);
    signal mulr_2_108 : std_logic_vector(9 downto 0);
    signal mulr_3_108 : std_logic_vector(9 downto 0);
    signal mulr_4_108 : std_logic_vector(9 downto 0);
    signal mulr_1_109 : std_logic_vector(9 downto 0);
    signal mulr_2_109 : std_logic_vector(9 downto 0);
    signal mulr_3_109 : std_logic_vector(9 downto 0);
    signal mulr_4_109 : std_logic_vector(9 downto 0);
    signal mulr_1_110 : std_logic_vector(9 downto 0);
    signal mulr_2_110 : std_logic_vector(9 downto 0);
    signal mulr_3_110 : std_logic_vector(9 downto 0);
    signal mulr_4_110 : std_logic_vector(9 downto 0);
    signal mulr_1_111 : std_logic_vector(9 downto 0);
    signal mulr_2_111 : std_logic_vector(9 downto 0);
    signal mulr_3_111 : std_logic_vector(9 downto 0);
    signal mulr_4_111 : std_logic_vector(9 downto 0);
    signal mulr_1_112 : std_logic_vector(9 downto 0);
    signal mulr_2_112 : std_logic_vector(9 downto 0);
    signal mulr_3_112 : std_logic_vector(9 downto 0);
    signal mulr_4_112 : std_logic_vector(9 downto 0);
    signal mulr_1_113 : std_logic_vector(9 downto 0);
    signal mulr_2_113 : std_logic_vector(9 downto 0);
    signal mulr_3_113 : std_logic_vector(9 downto 0);
    signal mulr_4_113 : std_logic_vector(9 downto 0);
    signal mulr_1_114 : std_logic_vector(9 downto 0);
    signal mulr_2_114 : std_logic_vector(9 downto 0);
    signal mulr_3_114 : std_logic_vector(9 downto 0);
    signal mulr_4_114 : std_logic_vector(9 downto 0);
    signal mulr_1_115 : std_logic_vector(9 downto 0);
    signal mulr_2_115 : std_logic_vector(9 downto 0);
    signal mulr_3_115 : std_logic_vector(9 downto 0);
    signal mulr_4_115 : std_logic_vector(9 downto 0);
    signal mulr_1_116 : std_logic_vector(9 downto 0);
    signal mulr_2_116 : std_logic_vector(9 downto 0);
    signal mulr_3_116 : std_logic_vector(9 downto 0);
    signal mulr_4_116 : std_logic_vector(9 downto 0);
    signal mulr_1_117 : std_logic_vector(9 downto 0);
    signal mulr_2_117 : std_logic_vector(9 downto 0);
    signal mulr_3_117 : std_logic_vector(9 downto 0);
    signal mulr_4_117 : std_logic_vector(9 downto 0);
    signal mulr_1_118 : std_logic_vector(9 downto 0);
    signal mulr_2_118 : std_logic_vector(9 downto 0);
    signal mulr_3_118 : std_logic_vector(9 downto 0);
    signal mulr_4_118 : std_logic_vector(9 downto 0);
    signal mulr_1_119 : std_logic_vector(9 downto 0);
    signal mulr_2_119 : std_logic_vector(9 downto 0);
    signal mulr_3_119 : std_logic_vector(9 downto 0);
    signal mulr_4_119 : std_logic_vector(9 downto 0);
    signal mulr_1_120 : std_logic_vector(9 downto 0);
    signal mulr_2_120 : std_logic_vector(9 downto 0);
    signal mulr_3_120 : std_logic_vector(9 downto 0);
    signal mulr_4_120 : std_logic_vector(9 downto 0);
    signal mulr_1_121 : std_logic_vector(9 downto 0);
    signal mulr_2_121 : std_logic_vector(9 downto 0);
    signal mulr_3_121 : std_logic_vector(9 downto 0);
    signal mulr_4_121 : std_logic_vector(9 downto 0);
    signal mulr_1_122 : std_logic_vector(9 downto 0);
    signal mulr_2_122 : std_logic_vector(9 downto 0);
    signal mulr_3_122 : std_logic_vector(9 downto 0);
    signal mulr_4_122 : std_logic_vector(9 downto 0);
    signal mulr_1_123 : std_logic_vector(9 downto 0);
    signal mulr_2_123 : std_logic_vector(9 downto 0);
    signal mulr_3_123 : std_logic_vector(9 downto 0);
    signal mulr_4_123 : std_logic_vector(9 downto 0);
    signal mulr_1_124 : std_logic_vector(9 downto 0);
    signal mulr_2_124 : std_logic_vector(9 downto 0);
    signal mulr_3_124 : std_logic_vector(9 downto 0);
    signal mulr_4_124 : std_logic_vector(9 downto 0);
    signal mulr_1_125 : std_logic_vector(9 downto 0);
    signal mulr_2_125 : std_logic_vector(9 downto 0);
    signal mulr_3_125 : std_logic_vector(9 downto 0);
    signal mulr_4_125 : std_logic_vector(9 downto 0);
    signal mulr_1_126 : std_logic_vector(9 downto 0);
    signal mulr_2_126 : std_logic_vector(9 downto 0);
    signal mulr_3_126 : std_logic_vector(9 downto 0);
    signal mulr_4_126 : std_logic_vector(9 downto 0);
    signal mulr_1_127 : std_logic_vector(9 downto 0);
    signal mulr_2_127 : std_logic_vector(9 downto 0);
    signal mulr_3_127 : std_logic_vector(9 downto 0);
    signal mulr_4_127 : std_logic_vector(9 downto 0);
    signal mulr_1_128 : std_logic_vector(9 downto 0);
    signal mulr_2_128 : std_logic_vector(9 downto 0);
    signal mulr_3_128 : std_logic_vector(9 downto 0);
    signal mulr_4_128 : std_logic_vector(9 downto 0);
    signal mulr_1_129 : std_logic_vector(9 downto 0);
    signal mulr_2_129 : std_logic_vector(9 downto 0);
    signal mulr_3_129 : std_logic_vector(9 downto 0);
    signal mulr_4_129 : std_logic_vector(9 downto 0);
    signal mulr_1_130 : std_logic_vector(9 downto 0);
    signal mulr_2_130 : std_logic_vector(9 downto 0);
    signal mulr_3_130 : std_logic_vector(9 downto 0);
    signal mulr_4_130 : std_logic_vector(9 downto 0);
    signal mulr_1_131 : std_logic_vector(9 downto 0);
    signal mulr_2_131 : std_logic_vector(9 downto 0);
    signal mulr_3_131 : std_logic_vector(9 downto 0);
    signal mulr_4_131 : std_logic_vector(9 downto 0);
    signal mulr_1_132 : std_logic_vector(9 downto 0);
    signal mulr_2_132 : std_logic_vector(9 downto 0);
    signal mulr_3_132 : std_logic_vector(9 downto 0);
    signal mulr_4_132 : std_logic_vector(9 downto 0);
    signal mulr_1_133 : std_logic_vector(9 downto 0);
    signal mulr_2_133 : std_logic_vector(9 downto 0);
    signal mulr_3_133 : std_logic_vector(9 downto 0);
    signal mulr_4_133 : std_logic_vector(9 downto 0);
    signal mulr_1_134 : std_logic_vector(9 downto 0);
    signal mulr_2_134 : std_logic_vector(9 downto 0);
    signal mulr_3_134 : std_logic_vector(9 downto 0);
    signal mulr_4_134 : std_logic_vector(9 downto 0);
    signal mulr_1_135 : std_logic_vector(9 downto 0);
    signal mulr_2_135 : std_logic_vector(9 downto 0);
    signal mulr_3_135 : std_logic_vector(9 downto 0);
    signal mulr_4_135 : std_logic_vector(9 downto 0);
    signal mulr_1_136 : std_logic_vector(9 downto 0);
    signal mulr_2_136 : std_logic_vector(9 downto 0);
    signal mulr_3_136 : std_logic_vector(9 downto 0);
    signal mulr_4_136 : std_logic_vector(9 downto 0);
    signal mulr_1_137 : std_logic_vector(9 downto 0);
    signal mulr_2_137 : std_logic_vector(9 downto 0);
    signal mulr_3_137 : std_logic_vector(9 downto 0);
    signal mulr_4_137 : std_logic_vector(9 downto 0);
    signal mulr_1_138 : std_logic_vector(9 downto 0);
    signal mulr_2_138 : std_logic_vector(9 downto 0);
    signal mulr_3_138 : std_logic_vector(9 downto 0);
    signal mulr_4_138 : std_logic_vector(9 downto 0);
    signal mulr_1_139 : std_logic_vector(9 downto 0);
    signal mulr_2_139 : std_logic_vector(9 downto 0);
    signal mulr_3_139 : std_logic_vector(9 downto 0);
    signal mulr_4_139 : std_logic_vector(9 downto 0);
    signal mulr_1_140 : std_logic_vector(9 downto 0);
    signal mulr_2_140 : std_logic_vector(9 downto 0);
    signal mulr_3_140 : std_logic_vector(9 downto 0);
    signal mulr_4_140 : std_logic_vector(9 downto 0);
    signal mulr_1_141 : std_logic_vector(9 downto 0);
    signal mulr_2_141 : std_logic_vector(9 downto 0);
    signal mulr_3_141 : std_logic_vector(9 downto 0);
    signal mulr_4_141 : std_logic_vector(9 downto 0);
    signal mulr_1_142 : std_logic_vector(9 downto 0);
    signal mulr_2_142 : std_logic_vector(9 downto 0);
    signal mulr_3_142 : std_logic_vector(9 downto 0);
    signal mulr_4_142 : std_logic_vector(9 downto 0);
    signal mulr_1_143 : std_logic_vector(9 downto 0);
    signal mulr_2_143 : std_logic_vector(9 downto 0);
    signal mulr_3_143 : std_logic_vector(9 downto 0);
    signal mulr_4_143 : std_logic_vector(9 downto 0);
    signal mulr_1_144 : std_logic_vector(9 downto 0);
    signal mulr_2_144 : std_logic_vector(9 downto 0);
    signal mulr_3_144 : std_logic_vector(9 downto 0);
    signal mulr_4_144 : std_logic_vector(9 downto 0);
    signal mulr_1_145 : std_logic_vector(9 downto 0);
    signal mulr_2_145 : std_logic_vector(9 downto 0);
    signal mulr_3_145 : std_logic_vector(9 downto 0);
    signal mulr_4_145 : std_logic_vector(9 downto 0);
    signal mulr_1_146 : std_logic_vector(9 downto 0);
    signal mulr_2_146 : std_logic_vector(9 downto 0);
    signal mulr_3_146 : std_logic_vector(9 downto 0);
    signal mulr_4_146 : std_logic_vector(9 downto 0);
    signal mulr_1_147 : std_logic_vector(9 downto 0);
    signal mulr_2_147 : std_logic_vector(9 downto 0);
    signal mulr_3_147 : std_logic_vector(9 downto 0);
    signal mulr_4_147 : std_logic_vector(9 downto 0);
    signal mulr_1_148 : std_logic_vector(9 downto 0);
    signal mulr_2_148 : std_logic_vector(9 downto 0);
    signal mulr_3_148 : std_logic_vector(9 downto 0);
    signal mulr_4_148 : std_logic_vector(9 downto 0);
    signal mulr_1_149 : std_logic_vector(9 downto 0);
    signal mulr_2_149 : std_logic_vector(9 downto 0);
    signal mulr_3_149 : std_logic_vector(9 downto 0);
    signal mulr_4_149 : std_logic_vector(9 downto 0);
    signal mulr_1_150 : std_logic_vector(9 downto 0);
    signal mulr_2_150 : std_logic_vector(9 downto 0);
    signal mulr_3_150 : std_logic_vector(9 downto 0);
    signal mulr_4_150 : std_logic_vector(9 downto 0);
    signal mulr_1_151 : std_logic_vector(9 downto 0);
    signal mulr_2_151 : std_logic_vector(9 downto 0);
    signal mulr_3_151 : std_logic_vector(9 downto 0);
    signal mulr_4_151 : std_logic_vector(9 downto 0);
    signal mulr_1_152 : std_logic_vector(9 downto 0);
    signal mulr_2_152 : std_logic_vector(9 downto 0);
    signal mulr_3_152 : std_logic_vector(9 downto 0);
    signal mulr_4_152 : std_logic_vector(9 downto 0);
    signal mulr_1_153 : std_logic_vector(9 downto 0);
    signal mulr_2_153 : std_logic_vector(9 downto 0);
    signal mulr_3_153 : std_logic_vector(9 downto 0);
    signal mulr_4_153 : std_logic_vector(9 downto 0);
    signal mulr_1_154 : std_logic_vector(9 downto 0);
    signal mulr_2_154 : std_logic_vector(9 downto 0);
    signal mulr_3_154 : std_logic_vector(9 downto 0);
    signal mulr_4_154 : std_logic_vector(9 downto 0);
    signal mulr_1_155 : std_logic_vector(9 downto 0);
    signal mulr_2_155 : std_logic_vector(9 downto 0);
    signal mulr_3_155 : std_logic_vector(9 downto 0);
    signal mulr_4_155 : std_logic_vector(9 downto 0);
    signal mulr_1_156 : std_logic_vector(9 downto 0);
    signal mulr_2_156 : std_logic_vector(9 downto 0);
    signal mulr_3_156 : std_logic_vector(9 downto 0);
    signal mulr_4_156 : std_logic_vector(9 downto 0);
    signal mulr_1_157 : std_logic_vector(9 downto 0);
    signal mulr_2_157 : std_logic_vector(9 downto 0);
    signal mulr_3_157 : std_logic_vector(9 downto 0);
    signal mulr_4_157 : std_logic_vector(9 downto 0);
    signal mulr_1_158 : std_logic_vector(9 downto 0);
    signal mulr_2_158 : std_logic_vector(9 downto 0);
    signal mulr_3_158 : std_logic_vector(9 downto 0);
    signal mulr_4_158 : std_logic_vector(9 downto 0);
    signal mulr_1_159 : std_logic_vector(9 downto 0);
    signal mulr_2_159 : std_logic_vector(9 downto 0);
    signal mulr_3_159 : std_logic_vector(9 downto 0);
    signal mulr_4_159 : std_logic_vector(9 downto 0);
    signal mulr_1_160 : std_logic_vector(9 downto 0);
    signal mulr_2_160 : std_logic_vector(9 downto 0);
    signal mulr_3_160 : std_logic_vector(9 downto 0);
    signal mulr_4_160 : std_logic_vector(9 downto 0);
    signal mulr_1_161 : std_logic_vector(9 downto 0);
    signal mulr_2_161 : std_logic_vector(9 downto 0);
    signal mulr_3_161 : std_logic_vector(9 downto 0);
    signal mulr_4_161 : std_logic_vector(9 downto 0);
    signal mulr_1_162 : std_logic_vector(9 downto 0);
    signal mulr_2_162 : std_logic_vector(9 downto 0);
    signal mulr_3_162 : std_logic_vector(9 downto 0);
    signal mulr_4_162 : std_logic_vector(9 downto 0);
    signal mulr_1_163 : std_logic_vector(9 downto 0);
    signal mulr_2_163 : std_logic_vector(9 downto 0);
    signal mulr_3_163 : std_logic_vector(9 downto 0);
    signal mulr_4_163 : std_logic_vector(9 downto 0);
    signal mulr_1_164 : std_logic_vector(9 downto 0);
    signal mulr_2_164 : std_logic_vector(9 downto 0);
    signal mulr_3_164 : std_logic_vector(9 downto 0);
    signal mulr_4_164 : std_logic_vector(9 downto 0);
    signal mulr_1_165 : std_logic_vector(9 downto 0);
    signal mulr_2_165 : std_logic_vector(9 downto 0);
    signal mulr_3_165 : std_logic_vector(9 downto 0);
    signal mulr_4_165 : std_logic_vector(9 downto 0);
    signal mulr_1_166 : std_logic_vector(9 downto 0);
    signal mulr_2_166 : std_logic_vector(9 downto 0);
    signal mulr_3_166 : std_logic_vector(9 downto 0);
    signal mulr_4_166 : std_logic_vector(9 downto 0);
    signal mulr_1_167 : std_logic_vector(9 downto 0);
    signal mulr_2_167 : std_logic_vector(9 downto 0);
    signal mulr_3_167 : std_logic_vector(9 downto 0);
    signal mulr_4_167 : std_logic_vector(9 downto 0);
    signal mulr_1_168 : std_logic_vector(9 downto 0);
    signal mulr_2_168 : std_logic_vector(9 downto 0);
    signal mulr_3_168 : std_logic_vector(9 downto 0);
    signal mulr_4_168 : std_logic_vector(9 downto 0);
    signal mulr_1_169 : std_logic_vector(9 downto 0);
    signal mulr_2_169 : std_logic_vector(9 downto 0);
    signal mulr_3_169 : std_logic_vector(9 downto 0);
    signal mulr_4_169 : std_logic_vector(9 downto 0);
    signal mulr_1_170 : std_logic_vector(9 downto 0);
    signal mulr_2_170 : std_logic_vector(9 downto 0);
    signal mulr_3_170 : std_logic_vector(9 downto 0);
    signal mulr_4_170 : std_logic_vector(9 downto 0);
    signal mulr_1_171 : std_logic_vector(9 downto 0);
    signal mulr_2_171 : std_logic_vector(9 downto 0);
    signal mulr_3_171 : std_logic_vector(9 downto 0);
    signal mulr_4_171 : std_logic_vector(9 downto 0);
    signal mulr_1_172 : std_logic_vector(9 downto 0);
    signal mulr_2_172 : std_logic_vector(9 downto 0);
    signal mulr_3_172 : std_logic_vector(9 downto 0);
    signal mulr_4_172 : std_logic_vector(9 downto 0);
    signal mulr_1_173 : std_logic_vector(9 downto 0);
    signal mulr_2_173 : std_logic_vector(9 downto 0);
    signal mulr_3_173 : std_logic_vector(9 downto 0);
    signal mulr_4_173 : std_logic_vector(9 downto 0);
    signal mulr_1_174 : std_logic_vector(9 downto 0);
    signal mulr_2_174 : std_logic_vector(9 downto 0);
    signal mulr_3_174 : std_logic_vector(9 downto 0);
    signal mulr_4_174 : std_logic_vector(9 downto 0);
    signal mulr_1_175 : std_logic_vector(9 downto 0);
    signal mulr_2_175 : std_logic_vector(9 downto 0);
    signal mulr_3_175 : std_logic_vector(9 downto 0);
    signal mulr_4_175 : std_logic_vector(9 downto 0);
    signal mulr_1_176 : std_logic_vector(9 downto 0);
    signal mulr_2_176 : std_logic_vector(9 downto 0);
    signal mulr_3_176 : std_logic_vector(9 downto 0);
    signal mulr_4_176 : std_logic_vector(9 downto 0);
    signal mulr_1_177 : std_logic_vector(9 downto 0);
    signal mulr_2_177 : std_logic_vector(9 downto 0);
    signal mulr_3_177 : std_logic_vector(9 downto 0);
    signal mulr_4_177 : std_logic_vector(9 downto 0);
    signal mulr_1_178 : std_logic_vector(9 downto 0);
    signal mulr_2_178 : std_logic_vector(9 downto 0);
    signal mulr_3_178 : std_logic_vector(9 downto 0);
    signal mulr_4_178 : std_logic_vector(9 downto 0);
    signal mulr_1_179 : std_logic_vector(9 downto 0);
    signal mulr_2_179 : std_logic_vector(9 downto 0);
    signal mulr_3_179 : std_logic_vector(9 downto 0);
    signal mulr_4_179 : std_logic_vector(9 downto 0);
    signal mulr_1_180 : std_logic_vector(9 downto 0);
    signal mulr_2_180 : std_logic_vector(9 downto 0);
    signal mulr_3_180 : std_logic_vector(9 downto 0);
    signal mulr_4_180 : std_logic_vector(9 downto 0);
    signal mulr_1_181 : std_logic_vector(9 downto 0);
    signal mulr_2_181 : std_logic_vector(9 downto 0);
    signal mulr_3_181 : std_logic_vector(9 downto 0);
    signal mulr_4_181 : std_logic_vector(9 downto 0);
    signal mulr_1_182 : std_logic_vector(9 downto 0);
    signal mulr_2_182 : std_logic_vector(9 downto 0);
    signal mulr_3_182 : std_logic_vector(9 downto 0);
    signal mulr_4_182 : std_logic_vector(9 downto 0);
    signal mulr_1_183 : std_logic_vector(9 downto 0);
    signal mulr_2_183 : std_logic_vector(9 downto 0);
    signal mulr_3_183 : std_logic_vector(9 downto 0);
    signal mulr_4_183 : std_logic_vector(9 downto 0);
    signal mulr_1_184 : std_logic_vector(9 downto 0);
    signal mulr_2_184 : std_logic_vector(9 downto 0);
    signal mulr_3_184 : std_logic_vector(9 downto 0);
    signal mulr_4_184 : std_logic_vector(9 downto 0);
    signal mulr_1_185 : std_logic_vector(9 downto 0);
    signal mulr_2_185 : std_logic_vector(9 downto 0);
    signal mulr_3_185 : std_logic_vector(9 downto 0);
    signal mulr_4_185 : std_logic_vector(9 downto 0);
    signal mulr_1_186 : std_logic_vector(9 downto 0);
    signal mulr_2_186 : std_logic_vector(9 downto 0);
    signal mulr_3_186 : std_logic_vector(9 downto 0);
    signal mulr_4_186 : std_logic_vector(9 downto 0);
    signal mulr_1_187 : std_logic_vector(9 downto 0);
    signal mulr_2_187 : std_logic_vector(9 downto 0);
    signal mulr_3_187 : std_logic_vector(9 downto 0);
    signal mulr_4_187 : std_logic_vector(9 downto 0);
    signal mulr_1_188 : std_logic_vector(9 downto 0);
    signal mulr_2_188 : std_logic_vector(9 downto 0);
    signal mulr_3_188 : std_logic_vector(9 downto 0);
    signal mulr_4_188 : std_logic_vector(9 downto 0);
    signal mulr_1_189 : std_logic_vector(9 downto 0);
    signal mulr_2_189 : std_logic_vector(9 downto 0);
    signal mulr_3_189 : std_logic_vector(9 downto 0);
    signal mulr_4_189 : std_logic_vector(9 downto 0);
    signal mulr_1_190 : std_logic_vector(9 downto 0);
    signal mulr_2_190 : std_logic_vector(9 downto 0);
    signal mulr_3_190 : std_logic_vector(9 downto 0);
    signal mulr_4_190 : std_logic_vector(9 downto 0);
    signal mulr_1_191 : std_logic_vector(9 downto 0);
    signal mulr_2_191 : std_logic_vector(9 downto 0);
    signal mulr_3_191 : std_logic_vector(9 downto 0);
    signal mulr_4_191 : std_logic_vector(9 downto 0);
    signal mulr_1_192 : std_logic_vector(9 downto 0);
    signal mulr_2_192 : std_logic_vector(9 downto 0);
    signal mulr_3_192 : std_logic_vector(9 downto 0);
    signal mulr_4_192 : std_logic_vector(9 downto 0);
    signal mulr_1_193 : std_logic_vector(9 downto 0);
    signal mulr_2_193 : std_logic_vector(9 downto 0);
    signal mulr_3_193 : std_logic_vector(9 downto 0);
    signal mulr_4_193 : std_logic_vector(9 downto 0);
    signal mulr_1_194 : std_logic_vector(9 downto 0);
    signal mulr_2_194 : std_logic_vector(9 downto 0);
    signal mulr_3_194 : std_logic_vector(9 downto 0);
    signal mulr_4_194 : std_logic_vector(9 downto 0);
    signal mulr_1_195 : std_logic_vector(9 downto 0);
    signal mulr_2_195 : std_logic_vector(9 downto 0);
    signal mulr_3_195 : std_logic_vector(9 downto 0);
    signal mulr_4_195 : std_logic_vector(9 downto 0);
    signal mulr_1_196 : std_logic_vector(9 downto 0);
    signal mulr_2_196 : std_logic_vector(9 downto 0);
    signal mulr_3_196 : std_logic_vector(9 downto 0);
    signal mulr_4_196 : std_logic_vector(9 downto 0);
    signal mulr_1_197 : std_logic_vector(9 downto 0);
    signal mulr_2_197 : std_logic_vector(9 downto 0);
    signal mulr_3_197 : std_logic_vector(9 downto 0);
    signal mulr_4_197 : std_logic_vector(9 downto 0);
    signal mulr_1_198 : std_logic_vector(9 downto 0);
    signal mulr_2_198 : std_logic_vector(9 downto 0);
    signal mulr_3_198 : std_logic_vector(9 downto 0);
    signal mulr_4_198 : std_logic_vector(9 downto 0);
    signal mulr_1_199 : std_logic_vector(9 downto 0);
    signal mulr_2_199 : std_logic_vector(9 downto 0);
    signal mulr_3_199 : std_logic_vector(9 downto 0);
    signal mulr_4_199 : std_logic_vector(9 downto 0);
    signal mulr_1_200 : std_logic_vector(9 downto 0);
    signal mulr_2_200 : std_logic_vector(9 downto 0);
    signal mulr_3_200 : std_logic_vector(9 downto 0);
    signal mulr_4_200 : std_logic_vector(9 downto 0);
    signal mulr_1_201 : std_logic_vector(9 downto 0);
    signal mulr_2_201 : std_logic_vector(9 downto 0);
    signal mulr_3_201 : std_logic_vector(9 downto 0);
    signal mulr_4_201 : std_logic_vector(9 downto 0);
    signal mulr_1_202 : std_logic_vector(9 downto 0);
    signal mulr_2_202 : std_logic_vector(9 downto 0);
    signal mulr_3_202 : std_logic_vector(9 downto 0);
    signal mulr_4_202 : std_logic_vector(9 downto 0);
    signal mulr_1_203 : std_logic_vector(9 downto 0);
    signal mulr_2_203 : std_logic_vector(9 downto 0);
    signal mulr_3_203 : std_logic_vector(9 downto 0);
    signal mulr_4_203 : std_logic_vector(9 downto 0);
    signal mulr_1_204 : std_logic_vector(9 downto 0);
    signal mulr_2_204 : std_logic_vector(9 downto 0);
    signal mulr_3_204 : std_logic_vector(9 downto 0);
    signal mulr_4_204 : std_logic_vector(9 downto 0);
    signal mulr_1_205 : std_logic_vector(9 downto 0);
    signal mulr_2_205 : std_logic_vector(9 downto 0);
    signal mulr_3_205 : std_logic_vector(9 downto 0);
    signal mulr_4_205 : std_logic_vector(9 downto 0);
    signal mulr_1_206 : std_logic_vector(9 downto 0);
    signal mulr_2_206 : std_logic_vector(9 downto 0);
    signal mulr_3_206 : std_logic_vector(9 downto 0);
    signal mulr_4_206 : std_logic_vector(9 downto 0);
    signal mulr_1_207 : std_logic_vector(9 downto 0);
    signal mulr_2_207 : std_logic_vector(9 downto 0);
    signal mulr_3_207 : std_logic_vector(9 downto 0);
    signal mulr_4_207 : std_logic_vector(9 downto 0);
    signal mulr_1_208 : std_logic_vector(9 downto 0);
    signal mulr_2_208 : std_logic_vector(9 downto 0);
    signal mulr_3_208 : std_logic_vector(9 downto 0);
    signal mulr_4_208 : std_logic_vector(9 downto 0);
    signal mulr_1_209 : std_logic_vector(9 downto 0);
    signal mulr_2_209 : std_logic_vector(9 downto 0);
    signal mulr_3_209 : std_logic_vector(9 downto 0);
    signal mulr_4_209 : std_logic_vector(9 downto 0);
    signal mulr_1_210 : std_logic_vector(9 downto 0);
    signal mulr_2_210 : std_logic_vector(9 downto 0);
    signal mulr_3_210 : std_logic_vector(9 downto 0);
    signal mulr_4_210 : std_logic_vector(9 downto 0);
    signal mulr_1_211 : std_logic_vector(9 downto 0);
    signal mulr_2_211 : std_logic_vector(9 downto 0);
    signal mulr_3_211 : std_logic_vector(9 downto 0);
    signal mulr_4_211 : std_logic_vector(9 downto 0);
    signal mulr_1_212 : std_logic_vector(9 downto 0);
    signal mulr_2_212 : std_logic_vector(9 downto 0);
    signal mulr_3_212 : std_logic_vector(9 downto 0);
    signal mulr_4_212 : std_logic_vector(9 downto 0);
    signal mulr_1_213 : std_logic_vector(9 downto 0);
    signal mulr_2_213 : std_logic_vector(9 downto 0);
    signal mulr_3_213 : std_logic_vector(9 downto 0);
    signal mulr_4_213 : std_logic_vector(9 downto 0);
    signal mulr_1_214 : std_logic_vector(9 downto 0);
    signal mulr_2_214 : std_logic_vector(9 downto 0);
    signal mulr_3_214 : std_logic_vector(9 downto 0);
    signal mulr_4_214 : std_logic_vector(9 downto 0);
    signal mulr_1_215 : std_logic_vector(9 downto 0);
    signal mulr_2_215 : std_logic_vector(9 downto 0);
    signal mulr_3_215 : std_logic_vector(9 downto 0);
    signal mulr_4_215 : std_logic_vector(9 downto 0);
    signal mulr_1_216 : std_logic_vector(9 downto 0);
    signal mulr_2_216 : std_logic_vector(9 downto 0);
    signal mulr_3_216 : std_logic_vector(9 downto 0);
    signal mulr_4_216 : std_logic_vector(9 downto 0);
    signal mulr_1_217 : std_logic_vector(9 downto 0);
    signal mulr_2_217 : std_logic_vector(9 downto 0);
    signal mulr_3_217 : std_logic_vector(9 downto 0);
    signal mulr_4_217 : std_logic_vector(9 downto 0);
    signal mulr_1_218 : std_logic_vector(9 downto 0);
    signal mulr_2_218 : std_logic_vector(9 downto 0);
    signal mulr_3_218 : std_logic_vector(9 downto 0);
    signal mulr_4_218 : std_logic_vector(9 downto 0);
    signal mulr_1_219 : std_logic_vector(9 downto 0);
    signal mulr_2_219 : std_logic_vector(9 downto 0);
    signal mulr_3_219 : std_logic_vector(9 downto 0);
    signal mulr_4_219 : std_logic_vector(9 downto 0);
    signal mulr_1_220 : std_logic_vector(9 downto 0);
    signal mulr_2_220 : std_logic_vector(9 downto 0);
    signal mulr_3_220 : std_logic_vector(9 downto 0);
    signal mulr_4_220 : std_logic_vector(9 downto 0);
    signal mulr_1_221 : std_logic_vector(9 downto 0);
    signal mulr_2_221 : std_logic_vector(9 downto 0);
    signal mulr_3_221 : std_logic_vector(9 downto 0);
    signal mulr_4_221 : std_logic_vector(9 downto 0);
    signal mulr_1_222 : std_logic_vector(9 downto 0);
    signal mulr_2_222 : std_logic_vector(9 downto 0);
    signal mulr_3_222 : std_logic_vector(9 downto 0);
    signal mulr_4_222 : std_logic_vector(9 downto 0);
    signal mulr_1_223 : std_logic_vector(9 downto 0);
    signal mulr_2_223 : std_logic_vector(9 downto 0);
    signal mulr_3_223 : std_logic_vector(9 downto 0);
    signal mulr_4_223 : std_logic_vector(9 downto 0);
    signal mulr_1_224 : std_logic_vector(9 downto 0);
    signal mulr_2_224 : std_logic_vector(9 downto 0);
    signal mulr_3_224 : std_logic_vector(9 downto 0);
    signal mulr_4_224 : std_logic_vector(9 downto 0);
    signal mulr_1_225 : std_logic_vector(9 downto 0);
    signal mulr_2_225 : std_logic_vector(9 downto 0);
    signal mulr_3_225 : std_logic_vector(9 downto 0);
    signal mulr_4_225 : std_logic_vector(9 downto 0);
    signal mulr_1_226 : std_logic_vector(9 downto 0);
    signal mulr_2_226 : std_logic_vector(9 downto 0);
    signal mulr_3_226 : std_logic_vector(9 downto 0);
    signal mulr_4_226 : std_logic_vector(9 downto 0);
    signal mulr_1_227 : std_logic_vector(9 downto 0);
    signal mulr_2_227 : std_logic_vector(9 downto 0);
    signal mulr_3_227 : std_logic_vector(9 downto 0);
    signal mulr_4_227 : std_logic_vector(9 downto 0);
    signal mulr_1_228 : std_logic_vector(9 downto 0);
    signal mulr_2_228 : std_logic_vector(9 downto 0);
    signal mulr_3_228 : std_logic_vector(9 downto 0);
    signal mulr_4_228 : std_logic_vector(9 downto 0);
    signal mulr_1_229 : std_logic_vector(9 downto 0);
    signal mulr_2_229 : std_logic_vector(9 downto 0);
    signal mulr_3_229 : std_logic_vector(9 downto 0);
    signal mulr_4_229 : std_logic_vector(9 downto 0);
    signal mulr_1_230 : std_logic_vector(9 downto 0);
    signal mulr_2_230 : std_logic_vector(9 downto 0);
    signal mulr_3_230 : std_logic_vector(9 downto 0);
    signal mulr_4_230 : std_logic_vector(9 downto 0);
    signal mulr_1_231 : std_logic_vector(9 downto 0);
    signal mulr_2_231 : std_logic_vector(9 downto 0);
    signal mulr_3_231 : std_logic_vector(9 downto 0);
    signal mulr_4_231 : std_logic_vector(9 downto 0);
    signal mulr_1_232 : std_logic_vector(9 downto 0);
    signal mulr_2_232 : std_logic_vector(9 downto 0);
    signal mulr_3_232 : std_logic_vector(9 downto 0);
    signal mulr_4_232 : std_logic_vector(9 downto 0);
    signal mulr_1_233 : std_logic_vector(9 downto 0);
    signal mulr_2_233 : std_logic_vector(9 downto 0);
    signal mulr_3_233 : std_logic_vector(9 downto 0);
    signal mulr_4_233 : std_logic_vector(9 downto 0);
    signal mulr_1_234 : std_logic_vector(9 downto 0);
    signal mulr_2_234 : std_logic_vector(9 downto 0);
    signal mulr_3_234 : std_logic_vector(9 downto 0);
    signal mulr_4_234 : std_logic_vector(9 downto 0);
    signal mulr_1_235 : std_logic_vector(9 downto 0);
    signal mulr_2_235 : std_logic_vector(9 downto 0);
    signal mulr_3_235 : std_logic_vector(9 downto 0);
    signal mulr_4_235 : std_logic_vector(9 downto 0);
    signal mulr_1_236 : std_logic_vector(9 downto 0);
    signal mulr_2_236 : std_logic_vector(9 downto 0);
    signal mulr_3_236 : std_logic_vector(9 downto 0);
    signal mulr_4_236 : std_logic_vector(9 downto 0);
    signal mulr_1_237 : std_logic_vector(9 downto 0);
    signal mulr_2_237 : std_logic_vector(9 downto 0);
    signal mulr_3_237 : std_logic_vector(9 downto 0);
    signal mulr_4_237 : std_logic_vector(9 downto 0);
    signal mulr_1_238 : std_logic_vector(9 downto 0);
    signal mulr_2_238 : std_logic_vector(9 downto 0);
    signal mulr_3_238 : std_logic_vector(9 downto 0);
    signal mulr_4_238 : std_logic_vector(9 downto 0);
    signal mulr_1_239 : std_logic_vector(9 downto 0);
    signal mulr_2_239 : std_logic_vector(9 downto 0);
    signal mulr_3_239 : std_logic_vector(9 downto 0);
    signal mulr_4_239 : std_logic_vector(9 downto 0);
    signal mulr_1_240 : std_logic_vector(9 downto 0);
    signal mulr_2_240 : std_logic_vector(9 downto 0);
    signal mulr_3_240 : std_logic_vector(9 downto 0);
    signal mulr_4_240 : std_logic_vector(9 downto 0);
    signal mulr_1_241 : std_logic_vector(9 downto 0);
    signal mulr_2_241 : std_logic_vector(9 downto 0);
    signal mulr_3_241 : std_logic_vector(9 downto 0);
    signal mulr_4_241 : std_logic_vector(9 downto 0);
    signal mulr_1_242 : std_logic_vector(9 downto 0);
    signal mulr_2_242 : std_logic_vector(9 downto 0);
    signal mulr_3_242 : std_logic_vector(9 downto 0);
    signal mulr_4_242 : std_logic_vector(9 downto 0);
    signal mulr_1_243 : std_logic_vector(9 downto 0);
    signal mulr_2_243 : std_logic_vector(9 downto 0);
    signal mulr_3_243 : std_logic_vector(9 downto 0);
    signal mulr_4_243 : std_logic_vector(9 downto 0);
    signal mulr_1_244 : std_logic_vector(9 downto 0);
    signal mulr_2_244 : std_logic_vector(9 downto 0);
    signal mulr_3_244 : std_logic_vector(9 downto 0);
    signal mulr_4_244 : std_logic_vector(9 downto 0);
    signal mulr_1_245 : std_logic_vector(9 downto 0);
    signal mulr_2_245 : std_logic_vector(9 downto 0);
    signal mulr_3_245 : std_logic_vector(9 downto 0);
    signal mulr_4_245 : std_logic_vector(9 downto 0);
    signal mulr_1_246 : std_logic_vector(9 downto 0);
    signal mulr_2_246 : std_logic_vector(9 downto 0);
    signal mulr_3_246 : std_logic_vector(9 downto 0);
    signal mulr_4_246 : std_logic_vector(9 downto 0);
    signal mulr_1_247 : std_logic_vector(9 downto 0);
    signal mulr_2_247 : std_logic_vector(9 downto 0);
    signal mulr_3_247 : std_logic_vector(9 downto 0);
    signal mulr_4_247 : std_logic_vector(9 downto 0);
    signal mulr_1_248 : std_logic_vector(9 downto 0);
    signal mulr_2_248 : std_logic_vector(9 downto 0);
    signal mulr_3_248 : std_logic_vector(9 downto 0);
    signal mulr_4_248 : std_logic_vector(9 downto 0);
    signal mulr_1_249 : std_logic_vector(9 downto 0);
    signal mulr_2_249 : std_logic_vector(9 downto 0);
    signal mulr_3_249 : std_logic_vector(9 downto 0);
    signal mulr_4_249 : std_logic_vector(9 downto 0);
    signal mulr_1_250 : std_logic_vector(9 downto 0);
    signal mulr_2_250 : std_logic_vector(9 downto 0);
    signal mulr_3_250 : std_logic_vector(9 downto 0);
    signal mulr_4_250 : std_logic_vector(9 downto 0);
    signal mulr_1_251 : std_logic_vector(9 downto 0);
    signal mulr_2_251 : std_logic_vector(9 downto 0);
    signal mulr_3_251 : std_logic_vector(9 downto 0);
    signal mulr_4_251 : std_logic_vector(9 downto 0);
    signal mulr_1_252 : std_logic_vector(9 downto 0);
    signal mulr_2_252 : std_logic_vector(9 downto 0);
    signal mulr_3_252 : std_logic_vector(9 downto 0);
    signal mulr_4_252 : std_logic_vector(9 downto 0);
    signal mulr_1_253 : std_logic_vector(9 downto 0);
    signal mulr_2_253 : std_logic_vector(9 downto 0);
    signal mulr_3_253 : std_logic_vector(9 downto 0);
    signal mulr_4_253 : std_logic_vector(9 downto 0);
    signal mulr_1_254 : std_logic_vector(9 downto 0);
    signal mulr_2_254 : std_logic_vector(9 downto 0);
    signal mulr_3_254 : std_logic_vector(9 downto 0);
    signal mulr_4_254 : std_logic_vector(9 downto 0);
    signal mulr_1_255 : std_logic_vector(9 downto 0);
    signal mulr_2_255 : std_logic_vector(9 downto 0);
    signal mulr_3_255 : std_logic_vector(9 downto 0);
    signal mulr_4_255 : std_logic_vector(9 downto 0);
    signal mulr_1_256 : std_logic_vector(9 downto 0);
    signal mulr_2_256 : std_logic_vector(9 downto 0);
    signal mulr_3_256 : std_logic_vector(9 downto 0);
    signal mulr_4_256 : std_logic_vector(9 downto 0);
    signal mulr_1_257 : std_logic_vector(9 downto 0);
    signal mulr_2_257 : std_logic_vector(9 downto 0);
    signal mulr_3_257 : std_logic_vector(9 downto 0);
    signal mulr_4_257 : std_logic_vector(9 downto 0);
    signal mulr_1_258 : std_logic_vector(9 downto 0);
    signal mulr_2_258 : std_logic_vector(9 downto 0);
    signal mulr_3_258 : std_logic_vector(9 downto 0);
    signal mulr_4_258 : std_logic_vector(9 downto 0);
    signal mulr_1_259 : std_logic_vector(9 downto 0);
    signal mulr_2_259 : std_logic_vector(9 downto 0);
    signal mulr_3_259 : std_logic_vector(9 downto 0);
    signal mulr_4_259 : std_logic_vector(9 downto 0);
    signal mulr_1_260 : std_logic_vector(9 downto 0);
    signal mulr_2_260 : std_logic_vector(9 downto 0);
    signal mulr_3_260 : std_logic_vector(9 downto 0);
    signal mulr_4_260 : std_logic_vector(9 downto 0);
    signal mulr_1_261 : std_logic_vector(9 downto 0);
    signal mulr_2_261 : std_logic_vector(9 downto 0);
    signal mulr_3_261 : std_logic_vector(9 downto 0);
    signal mulr_4_261 : std_logic_vector(9 downto 0);
    signal mulr_1_262 : std_logic_vector(9 downto 0);
    signal mulr_2_262 : std_logic_vector(9 downto 0);
    signal mulr_3_262 : std_logic_vector(9 downto 0);
    signal mulr_4_262 : std_logic_vector(9 downto 0);
    signal mulr_1_263 : std_logic_vector(9 downto 0);
    signal mulr_2_263 : std_logic_vector(9 downto 0);
    signal mulr_3_263 : std_logic_vector(9 downto 0);
    signal mulr_4_263 : std_logic_vector(9 downto 0);
    signal mulr_1_264 : std_logic_vector(9 downto 0);
    signal mulr_2_264 : std_logic_vector(9 downto 0);
    signal mulr_3_264 : std_logic_vector(9 downto 0);
    signal mulr_4_264 : std_logic_vector(9 downto 0);
    signal mulr_1_265 : std_logic_vector(9 downto 0);
    signal mulr_2_265 : std_logic_vector(9 downto 0);
    signal mulr_3_265 : std_logic_vector(9 downto 0);
    signal mulr_4_265 : std_logic_vector(9 downto 0);
    signal mulr_1_266 : std_logic_vector(9 downto 0);
    signal mulr_2_266 : std_logic_vector(9 downto 0);
    signal mulr_3_266 : std_logic_vector(9 downto 0);
    signal mulr_4_266 : std_logic_vector(9 downto 0);
    signal mulr_1_267 : std_logic_vector(9 downto 0);
    signal mulr_2_267 : std_logic_vector(9 downto 0);
    signal mulr_3_267 : std_logic_vector(9 downto 0);
    signal mulr_4_267 : std_logic_vector(9 downto 0);
    signal mulr_1_268 : std_logic_vector(9 downto 0);
    signal mulr_2_268 : std_logic_vector(9 downto 0);
    signal mulr_3_268 : std_logic_vector(9 downto 0);
    signal mulr_4_268 : std_logic_vector(9 downto 0);
    signal mulr_1_269 : std_logic_vector(9 downto 0);
    signal mulr_2_269 : std_logic_vector(9 downto 0);
    signal mulr_3_269 : std_logic_vector(9 downto 0);
    signal mulr_4_269 : std_logic_vector(9 downto 0);
    signal mulr_1_270 : std_logic_vector(9 downto 0);
    signal mulr_2_270 : std_logic_vector(9 downto 0);
    signal mulr_3_270 : std_logic_vector(9 downto 0);
    signal mulr_4_270 : std_logic_vector(9 downto 0);
    signal mulr_1_271 : std_logic_vector(9 downto 0);
    signal mulr_2_271 : std_logic_vector(9 downto 0);
    signal mulr_3_271 : std_logic_vector(9 downto 0);
    signal mulr_4_271 : std_logic_vector(9 downto 0);
    signal mulr_1_272 : std_logic_vector(9 downto 0);
    signal mulr_2_272 : std_logic_vector(9 downto 0);
    signal mulr_3_272 : std_logic_vector(9 downto 0);
    signal mulr_4_272 : std_logic_vector(9 downto 0);
    signal mulr_1_273 : std_logic_vector(9 downto 0);
    signal mulr_2_273 : std_logic_vector(9 downto 0);
    signal mulr_3_273 : std_logic_vector(9 downto 0);
    signal mulr_4_273 : std_logic_vector(9 downto 0);
    signal mulr_1_274 : std_logic_vector(9 downto 0);
    signal mulr_2_274 : std_logic_vector(9 downto 0);
    signal mulr_3_274 : std_logic_vector(9 downto 0);
    signal mulr_4_274 : std_logic_vector(9 downto 0);
    signal mulr_1_275 : std_logic_vector(9 downto 0);
    signal mulr_2_275 : std_logic_vector(9 downto 0);
    signal mulr_3_275 : std_logic_vector(9 downto 0);
    signal mulr_4_275 : std_logic_vector(9 downto 0);
    signal mulr_1_276 : std_logic_vector(9 downto 0);
    signal mulr_2_276 : std_logic_vector(9 downto 0);
    signal mulr_3_276 : std_logic_vector(9 downto 0);
    signal mulr_4_276 : std_logic_vector(9 downto 0);
    signal mulr_1_277 : std_logic_vector(9 downto 0);
    signal mulr_2_277 : std_logic_vector(9 downto 0);
    signal mulr_3_277 : std_logic_vector(9 downto 0);
    signal mulr_4_277 : std_logic_vector(9 downto 0);
    signal mulr_1_278 : std_logic_vector(9 downto 0);
    signal mulr_2_278 : std_logic_vector(9 downto 0);
    signal mulr_3_278 : std_logic_vector(9 downto 0);
    signal mulr_4_278 : std_logic_vector(9 downto 0);
    signal mulr_1_279 : std_logic_vector(9 downto 0);
    signal mulr_2_279 : std_logic_vector(9 downto 0);
    signal mulr_3_279 : std_logic_vector(9 downto 0);
    signal mulr_4_279 : std_logic_vector(9 downto 0);
    signal mulr_1_280 : std_logic_vector(9 downto 0);
    signal mulr_2_280 : std_logic_vector(9 downto 0);
    signal mulr_3_280 : std_logic_vector(9 downto 0);
    signal mulr_4_280 : std_logic_vector(9 downto 0);
    signal mulr_1_281 : std_logic_vector(9 downto 0);
    signal mulr_2_281 : std_logic_vector(9 downto 0);
    signal mulr_3_281 : std_logic_vector(9 downto 0);
    signal mulr_4_281 : std_logic_vector(9 downto 0);
    signal mulr_1_282 : std_logic_vector(9 downto 0);
    signal mulr_2_282 : std_logic_vector(9 downto 0);
    signal mulr_3_282 : std_logic_vector(9 downto 0);
    signal mulr_4_282 : std_logic_vector(9 downto 0);
    signal mulr_1_283 : std_logic_vector(9 downto 0);
    signal mulr_2_283 : std_logic_vector(9 downto 0);
    signal mulr_3_283 : std_logic_vector(9 downto 0);
    signal mulr_4_283 : std_logic_vector(9 downto 0);
    signal mulr_1_284 : std_logic_vector(9 downto 0);
    signal mulr_2_284 : std_logic_vector(9 downto 0);
    signal mulr_3_284 : std_logic_vector(9 downto 0);
    signal mulr_4_284 : std_logic_vector(9 downto 0);
    signal mulr_1_285 : std_logic_vector(9 downto 0);
    signal mulr_2_285 : std_logic_vector(9 downto 0);
    signal mulr_3_285 : std_logic_vector(9 downto 0);
    signal mulr_4_285 : std_logic_vector(9 downto 0);
    signal mulr_1_286 : std_logic_vector(9 downto 0);
    signal mulr_2_286 : std_logic_vector(9 downto 0);
    signal mulr_3_286 : std_logic_vector(9 downto 0);
    signal mulr_4_286 : std_logic_vector(9 downto 0);
    signal mulr_1_287 : std_logic_vector(9 downto 0);
    signal mulr_2_287 : std_logic_vector(9 downto 0);
    signal mulr_3_287 : std_logic_vector(9 downto 0);
    signal mulr_4_287 : std_logic_vector(9 downto 0);
    signal mulr_1_288 : std_logic_vector(9 downto 0);
    signal mulr_2_288 : std_logic_vector(9 downto 0);
    signal mulr_3_288 : std_logic_vector(9 downto 0);
    signal mulr_4_288 : std_logic_vector(9 downto 0);
    signal mulr_1_289 : std_logic_vector(9 downto 0);
    signal mulr_2_289 : std_logic_vector(9 downto 0);
    signal mulr_3_289 : std_logic_vector(9 downto 0);
    signal mulr_4_289 : std_logic_vector(9 downto 0);
    signal mulr_1_290 : std_logic_vector(9 downto 0);
    signal mulr_2_290 : std_logic_vector(9 downto 0);
    signal mulr_3_290 : std_logic_vector(9 downto 0);
    signal mulr_4_290 : std_logic_vector(9 downto 0);
    signal mulr_1_291 : std_logic_vector(9 downto 0);
    signal mulr_2_291 : std_logic_vector(9 downto 0);
    signal mulr_3_291 : std_logic_vector(9 downto 0);
    signal mulr_4_291 : std_logic_vector(9 downto 0);
    signal mulr_1_292 : std_logic_vector(9 downto 0);
    signal mulr_2_292 : std_logic_vector(9 downto 0);
    signal mulr_3_292 : std_logic_vector(9 downto 0);
    signal mulr_4_292 : std_logic_vector(9 downto 0);
    signal mulr_1_293 : std_logic_vector(9 downto 0);
    signal mulr_2_293 : std_logic_vector(9 downto 0);
    signal mulr_3_293 : std_logic_vector(9 downto 0);
    signal mulr_4_293 : std_logic_vector(9 downto 0);
    signal mulr_1_294 : std_logic_vector(9 downto 0);
    signal mulr_2_294 : std_logic_vector(9 downto 0);
    signal mulr_3_294 : std_logic_vector(9 downto 0);
    signal mulr_4_294 : std_logic_vector(9 downto 0);
    signal mulr_1_295 : std_logic_vector(9 downto 0);
    signal mulr_2_295 : std_logic_vector(9 downto 0);
    signal mulr_3_295 : std_logic_vector(9 downto 0);
    signal mulr_4_295 : std_logic_vector(9 downto 0);
    signal mulr_1_296 : std_logic_vector(9 downto 0);
    signal mulr_2_296 : std_logic_vector(9 downto 0);
    signal mulr_3_296 : std_logic_vector(9 downto 0);
    signal mulr_4_296 : std_logic_vector(9 downto 0);
    signal mulr_1_297 : std_logic_vector(9 downto 0);
    signal mulr_2_297 : std_logic_vector(9 downto 0);
    signal mulr_3_297 : std_logic_vector(9 downto 0);
    signal mulr_4_297 : std_logic_vector(9 downto 0);
    signal mulr_1_298 : std_logic_vector(9 downto 0);
    signal mulr_2_298 : std_logic_vector(9 downto 0);
    signal mulr_3_298 : std_logic_vector(9 downto 0);
    signal mulr_4_298 : std_logic_vector(9 downto 0);
    signal mulr_1_299 : std_logic_vector(9 downto 0);
    signal mulr_2_299 : std_logic_vector(9 downto 0);
    signal mulr_3_299 : std_logic_vector(9 downto 0);
    signal mulr_4_299 : std_logic_vector(9 downto 0);
    signal mulr_1_300 : std_logic_vector(9 downto 0);
    signal mulr_2_300 : std_logic_vector(9 downto 0);
    signal mulr_3_300 : std_logic_vector(9 downto 0);
    signal mulr_4_300 : std_logic_vector(9 downto 0);
    signal mulr_1_301 : std_logic_vector(9 downto 0);
    signal mulr_2_301 : std_logic_vector(9 downto 0);
    signal mulr_3_301 : std_logic_vector(9 downto 0);
    signal mulr_4_301 : std_logic_vector(9 downto 0);
    signal mulr_1_302 : std_logic_vector(9 downto 0);
    signal mulr_2_302 : std_logic_vector(9 downto 0);
    signal mulr_3_302 : std_logic_vector(9 downto 0);
    signal mulr_4_302 : std_logic_vector(9 downto 0);
    signal mulr_1_303 : std_logic_vector(9 downto 0);
    signal mulr_2_303 : std_logic_vector(9 downto 0);
    signal mulr_3_303 : std_logic_vector(9 downto 0);
    signal mulr_4_303 : std_logic_vector(9 downto 0);
    signal mulr_1_304 : std_logic_vector(9 downto 0);
    signal mulr_2_304 : std_logic_vector(9 downto 0);
    signal mulr_3_304 : std_logic_vector(9 downto 0);
    signal mulr_4_304 : std_logic_vector(9 downto 0);
    signal mulr_1_305 : std_logic_vector(9 downto 0);
    signal mulr_2_305 : std_logic_vector(9 downto 0);
    signal mulr_3_305 : std_logic_vector(9 downto 0);
    signal mulr_4_305 : std_logic_vector(9 downto 0);
    signal mulr_1_306 : std_logic_vector(9 downto 0);
    signal mulr_2_306 : std_logic_vector(9 downto 0);
    signal mulr_3_306 : std_logic_vector(9 downto 0);
    signal mulr_4_306 : std_logic_vector(9 downto 0);
    signal mulr_1_307 : std_logic_vector(9 downto 0);
    signal mulr_2_307 : std_logic_vector(9 downto 0);
    signal mulr_3_307 : std_logic_vector(9 downto 0);
    signal mulr_4_307 : std_logic_vector(9 downto 0);
    signal mulr_1_308 : std_logic_vector(9 downto 0);
    signal mulr_2_308 : std_logic_vector(9 downto 0);
    signal mulr_3_308 : std_logic_vector(9 downto 0);
    signal mulr_4_308 : std_logic_vector(9 downto 0);
    signal mulr_1_309 : std_logic_vector(9 downto 0);
    signal mulr_2_309 : std_logic_vector(9 downto 0);
    signal mulr_3_309 : std_logic_vector(9 downto 0);
    signal mulr_4_309 : std_logic_vector(9 downto 0);
    signal mulr_1_310 : std_logic_vector(9 downto 0);
    signal mulr_2_310 : std_logic_vector(9 downto 0);
    signal mulr_3_310 : std_logic_vector(9 downto 0);
    signal mulr_4_310 : std_logic_vector(9 downto 0);
    signal mulr_1_311 : std_logic_vector(9 downto 0);
    signal mulr_2_311 : std_logic_vector(9 downto 0);
    signal mulr_3_311 : std_logic_vector(9 downto 0);
    signal mulr_4_311 : std_logic_vector(9 downto 0);
    signal mulr_1_312 : std_logic_vector(9 downto 0);
    signal mulr_2_312 : std_logic_vector(9 downto 0);
    signal mulr_3_312 : std_logic_vector(9 downto 0);
    signal mulr_4_312 : std_logic_vector(9 downto 0);
    signal mulr_1_313 : std_logic_vector(9 downto 0);
    signal mulr_2_313 : std_logic_vector(9 downto 0);
    signal mulr_3_313 : std_logic_vector(9 downto 0);
    signal mulr_4_313 : std_logic_vector(9 downto 0);
    signal mulr_1_314 : std_logic_vector(9 downto 0);
    signal mulr_2_314 : std_logic_vector(9 downto 0);
    signal mulr_3_314 : std_logic_vector(9 downto 0);
    signal mulr_4_314 : std_logic_vector(9 downto 0);
    signal mulr_1_315 : std_logic_vector(9 downto 0);
    signal mulr_2_315 : std_logic_vector(9 downto 0);
    signal mulr_3_315 : std_logic_vector(9 downto 0);
    signal mulr_4_315 : std_logic_vector(9 downto 0);
    signal mulr_1_316 : std_logic_vector(9 downto 0);
    signal mulr_2_316 : std_logic_vector(9 downto 0);
    signal mulr_3_316 : std_logic_vector(9 downto 0);
    signal mulr_4_316 : std_logic_vector(9 downto 0);
    signal mulr_1_317 : std_logic_vector(9 downto 0);
    signal mulr_2_317 : std_logic_vector(9 downto 0);
    signal mulr_3_317 : std_logic_vector(9 downto 0);
    signal mulr_4_317 : std_logic_vector(9 downto 0);
    signal mulr_1_318 : std_logic_vector(9 downto 0);
    signal mulr_2_318 : std_logic_vector(9 downto 0);
    signal mulr_3_318 : std_logic_vector(9 downto 0);
    signal mulr_4_318 : std_logic_vector(9 downto 0);
    signal mulr_1_319 : std_logic_vector(9 downto 0);
    signal mulr_2_319 : std_logic_vector(9 downto 0);
    signal mulr_3_319 : std_logic_vector(9 downto 0);
    signal mulr_4_319 : std_logic_vector(9 downto 0);
    signal mulr_1_320 : std_logic_vector(9 downto 0);
    signal mulr_2_320 : std_logic_vector(9 downto 0);
    signal mulr_3_320 : std_logic_vector(9 downto 0);
    signal mulr_4_320 : std_logic_vector(9 downto 0);
    signal mulr_1_321 : std_logic_vector(9 downto 0);
    signal mulr_2_321 : std_logic_vector(9 downto 0);
    signal mulr_3_321 : std_logic_vector(9 downto 0);
    signal mulr_4_321 : std_logic_vector(9 downto 0);
    signal mulr_1_322 : std_logic_vector(9 downto 0);
    signal mulr_2_322 : std_logic_vector(9 downto 0);
    signal mulr_3_322 : std_logic_vector(9 downto 0);
    signal mulr_4_322 : std_logic_vector(9 downto 0);
    signal mulr_1_323 : std_logic_vector(9 downto 0);
    signal mulr_2_323 : std_logic_vector(9 downto 0);
    signal mulr_3_323 : std_logic_vector(9 downto 0);
    signal mulr_4_323 : std_logic_vector(9 downto 0);
    signal mulr_1_324 : std_logic_vector(9 downto 0);
    signal mulr_2_324 : std_logic_vector(9 downto 0);
    signal mulr_3_324 : std_logic_vector(9 downto 0);
    signal mulr_4_324 : std_logic_vector(9 downto 0);
    signal mulr_1_325 : std_logic_vector(9 downto 0);
    signal mulr_2_325 : std_logic_vector(9 downto 0);
    signal mulr_3_325 : std_logic_vector(9 downto 0);
    signal mulr_4_325 : std_logic_vector(9 downto 0);
    signal mulr_1_326 : std_logic_vector(9 downto 0);
    signal mulr_2_326 : std_logic_vector(9 downto 0);
    signal mulr_3_326 : std_logic_vector(9 downto 0);
    signal mulr_4_326 : std_logic_vector(9 downto 0);
    signal mulr_1_327 : std_logic_vector(9 downto 0);
    signal mulr_2_327 : std_logic_vector(9 downto 0);
    signal mulr_3_327 : std_logic_vector(9 downto 0);
    signal mulr_4_327 : std_logic_vector(9 downto 0);
    signal mulr_1_328 : std_logic_vector(9 downto 0);
    signal mulr_2_328 : std_logic_vector(9 downto 0);
    signal mulr_3_328 : std_logic_vector(9 downto 0);
    signal mulr_4_328 : std_logic_vector(9 downto 0);
    signal mulr_1_329 : std_logic_vector(9 downto 0);
    signal mulr_2_329 : std_logic_vector(9 downto 0);
    signal mulr_3_329 : std_logic_vector(9 downto 0);
    signal mulr_4_329 : std_logic_vector(9 downto 0);
    signal mulr_1_330 : std_logic_vector(9 downto 0);
    signal mulr_2_330 : std_logic_vector(9 downto 0);
    signal mulr_3_330 : std_logic_vector(9 downto 0);
    signal mulr_4_330 : std_logic_vector(9 downto 0);
    signal mulr_1_331 : std_logic_vector(9 downto 0);
    signal mulr_2_331 : std_logic_vector(9 downto 0);
    signal mulr_3_331 : std_logic_vector(9 downto 0);
    signal mulr_4_331 : std_logic_vector(9 downto 0);
    signal mulr_1_332 : std_logic_vector(9 downto 0);
    signal mulr_2_332 : std_logic_vector(9 downto 0);
    signal mulr_3_332 : std_logic_vector(9 downto 0);
    signal mulr_4_332 : std_logic_vector(9 downto 0);
    signal mulr_1_333 : std_logic_vector(9 downto 0);
    signal mulr_2_333 : std_logic_vector(9 downto 0);
    signal mulr_3_333 : std_logic_vector(9 downto 0);
    signal mulr_4_333 : std_logic_vector(9 downto 0);
    signal mulr_1_334 : std_logic_vector(9 downto 0);
    signal mulr_2_334 : std_logic_vector(9 downto 0);
    signal mulr_3_334 : std_logic_vector(9 downto 0);
    signal mulr_4_334 : std_logic_vector(9 downto 0);
    signal mulr_1_335 : std_logic_vector(9 downto 0);
    signal mulr_2_335 : std_logic_vector(9 downto 0);
    signal mulr_3_335 : std_logic_vector(9 downto 0);
    signal mulr_4_335 : std_logic_vector(9 downto 0);
    signal mulr_1_336 : std_logic_vector(9 downto 0);
    signal mulr_2_336 : std_logic_vector(9 downto 0);
    signal mulr_3_336 : std_logic_vector(9 downto 0);
    signal mulr_4_336 : std_logic_vector(9 downto 0);
    signal mulr_1_337 : std_logic_vector(9 downto 0);
    signal mulr_2_337 : std_logic_vector(9 downto 0);
    signal mulr_3_337 : std_logic_vector(9 downto 0);
    signal mulr_4_337 : std_logic_vector(9 downto 0);
    signal mulr_1_338 : std_logic_vector(9 downto 0);
    signal mulr_2_338 : std_logic_vector(9 downto 0);
    signal mulr_3_338 : std_logic_vector(9 downto 0);
    signal mulr_4_338 : std_logic_vector(9 downto 0);
    signal mulr_1_339 : std_logic_vector(9 downto 0);
    signal mulr_2_339 : std_logic_vector(9 downto 0);
    signal mulr_3_339 : std_logic_vector(9 downto 0);
    signal mulr_4_339 : std_logic_vector(9 downto 0);
    signal mulr_1_340 : std_logic_vector(9 downto 0);
    signal mulr_2_340 : std_logic_vector(9 downto 0);
    signal mulr_3_340 : std_logic_vector(9 downto 0);
    signal mulr_4_340 : std_logic_vector(9 downto 0);
    signal mulr_1_341 : std_logic_vector(9 downto 0);
    signal mulr_2_341 : std_logic_vector(9 downto 0);
    signal mulr_3_341 : std_logic_vector(9 downto 0);
    signal mulr_4_341 : std_logic_vector(9 downto 0);
    signal mulr_1_342 : std_logic_vector(9 downto 0);
    signal mulr_2_342 : std_logic_vector(9 downto 0);
    signal mulr_3_342 : std_logic_vector(9 downto 0);
    signal mulr_4_342 : std_logic_vector(9 downto 0);
    signal mulr_1_343 : std_logic_vector(9 downto 0);
    signal mulr_2_343 : std_logic_vector(9 downto 0);
    signal mulr_3_343 : std_logic_vector(9 downto 0);
    signal mulr_4_343 : std_logic_vector(9 downto 0);
    signal mulr_1_344 : std_logic_vector(9 downto 0);
    signal mulr_2_344 : std_logic_vector(9 downto 0);
    signal mulr_3_344 : std_logic_vector(9 downto 0);
    signal mulr_4_344 : std_logic_vector(9 downto 0);
    signal mulr_1_345 : std_logic_vector(9 downto 0);
    signal mulr_2_345 : std_logic_vector(9 downto 0);
    signal mulr_3_345 : std_logic_vector(9 downto 0);
    signal mulr_4_345 : std_logic_vector(9 downto 0);
    signal mulr_1_346 : std_logic_vector(9 downto 0);
    signal mulr_2_346 : std_logic_vector(9 downto 0);
    signal mulr_3_346 : std_logic_vector(9 downto 0);
    signal mulr_4_346 : std_logic_vector(9 downto 0);
    signal mulr_1_347 : std_logic_vector(9 downto 0);
    signal mulr_2_347 : std_logic_vector(9 downto 0);
    signal mulr_3_347 : std_logic_vector(9 downto 0);
    signal mulr_4_347 : std_logic_vector(9 downto 0);
    signal mulr_1_348 : std_logic_vector(9 downto 0);
    signal mulr_2_348 : std_logic_vector(9 downto 0);
    signal mulr_3_348 : std_logic_vector(9 downto 0);
    signal mulr_4_348 : std_logic_vector(9 downto 0);
    signal mulr_1_349 : std_logic_vector(9 downto 0);
    signal mulr_2_349 : std_logic_vector(9 downto 0);
    signal mulr_3_349 : std_logic_vector(9 downto 0);
    signal mulr_4_349 : std_logic_vector(9 downto 0);
    signal mulr_1_350 : std_logic_vector(9 downto 0);
    signal mulr_2_350 : std_logic_vector(9 downto 0);
    signal mulr_3_350 : std_logic_vector(9 downto 0);
    signal mulr_4_350 : std_logic_vector(9 downto 0);
    signal mulr_1_351 : std_logic_vector(9 downto 0);
    signal mulr_2_351 : std_logic_vector(9 downto 0);
    signal mulr_3_351 : std_logic_vector(9 downto 0);
    signal mulr_4_351 : std_logic_vector(9 downto 0);
    signal mulr_1_352 : std_logic_vector(9 downto 0);
    signal mulr_2_352 : std_logic_vector(9 downto 0);
    signal mulr_3_352 : std_logic_vector(9 downto 0);
    signal mulr_4_352 : std_logic_vector(9 downto 0);
    signal mulr_1_353 : std_logic_vector(9 downto 0);
    signal mulr_2_353 : std_logic_vector(9 downto 0);
    signal mulr_3_353 : std_logic_vector(9 downto 0);
    signal mulr_4_353 : std_logic_vector(9 downto 0);
    signal mulr_1_354 : std_logic_vector(9 downto 0);
    signal mulr_2_354 : std_logic_vector(9 downto 0);
    signal mulr_3_354 : std_logic_vector(9 downto 0);
    signal mulr_4_354 : std_logic_vector(9 downto 0);
    signal mulr_1_355 : std_logic_vector(9 downto 0);
    signal mulr_2_355 : std_logic_vector(9 downto 0);
    signal mulr_3_355 : std_logic_vector(9 downto 0);
    signal mulr_4_355 : std_logic_vector(9 downto 0);
    signal mulr_1_356 : std_logic_vector(9 downto 0);
    signal mulr_2_356 : std_logic_vector(9 downto 0);
    signal mulr_3_356 : std_logic_vector(9 downto 0);
    signal mulr_4_356 : std_logic_vector(9 downto 0);
    signal mulr_1_357 : std_logic_vector(9 downto 0);
    signal mulr_2_357 : std_logic_vector(9 downto 0);
    signal mulr_3_357 : std_logic_vector(9 downto 0);
    signal mulr_4_357 : std_logic_vector(9 downto 0);
    signal mulr_1_358 : std_logic_vector(9 downto 0);
    signal mulr_2_358 : std_logic_vector(9 downto 0);
    signal mulr_3_358 : std_logic_vector(9 downto 0);
    signal mulr_4_358 : std_logic_vector(9 downto 0);
    signal mulr_1_359 : std_logic_vector(9 downto 0);
    signal mulr_2_359 : std_logic_vector(9 downto 0);
    signal mulr_3_359 : std_logic_vector(9 downto 0);
    signal mulr_4_359 : std_logic_vector(9 downto 0);
    signal mulr_1_360 : std_logic_vector(9 downto 0);
    signal mulr_2_360 : std_logic_vector(9 downto 0);
    signal mulr_3_360 : std_logic_vector(9 downto 0);
    signal mulr_4_360 : std_logic_vector(9 downto 0);
    signal mulr_1_361 : std_logic_vector(9 downto 0);
    signal mulr_2_361 : std_logic_vector(9 downto 0);
    signal mulr_3_361 : std_logic_vector(9 downto 0);
    signal mulr_4_361 : std_logic_vector(9 downto 0);
    signal mulr_1_362 : std_logic_vector(9 downto 0);
    signal mulr_2_362 : std_logic_vector(9 downto 0);
    signal mulr_3_362 : std_logic_vector(9 downto 0);
    signal mulr_4_362 : std_logic_vector(9 downto 0);
    signal mulr_1_363 : std_logic_vector(9 downto 0);
    signal mulr_2_363 : std_logic_vector(9 downto 0);
    signal mulr_3_363 : std_logic_vector(9 downto 0);
    signal mulr_4_363 : std_logic_vector(9 downto 0);
    signal mulr_1_364 : std_logic_vector(9 downto 0);
    signal mulr_2_364 : std_logic_vector(9 downto 0);
    signal mulr_3_364 : std_logic_vector(9 downto 0);
    signal mulr_4_364 : std_logic_vector(9 downto 0);
    signal mulr_1_365 : std_logic_vector(9 downto 0);
    signal mulr_2_365 : std_logic_vector(9 downto 0);
    signal mulr_3_365 : std_logic_vector(9 downto 0);
    signal mulr_4_365 : std_logic_vector(9 downto 0);
    signal mulr_1_366 : std_logic_vector(9 downto 0);
    signal mulr_2_366 : std_logic_vector(9 downto 0);
    signal mulr_3_366 : std_logic_vector(9 downto 0);
    signal mulr_4_366 : std_logic_vector(9 downto 0);
    signal mulr_1_367 : std_logic_vector(9 downto 0);
    signal mulr_2_367 : std_logic_vector(9 downto 0);
    signal mulr_3_367 : std_logic_vector(9 downto 0);
    signal mulr_4_367 : std_logic_vector(9 downto 0);
    signal mulr_1_368 : std_logic_vector(9 downto 0);
    signal mulr_2_368 : std_logic_vector(9 downto 0);
    signal mulr_3_368 : std_logic_vector(9 downto 0);
    signal mulr_4_368 : std_logic_vector(9 downto 0);
    signal mulr_1_369 : std_logic_vector(9 downto 0);
    signal mulr_2_369 : std_logic_vector(9 downto 0);
    signal mulr_3_369 : std_logic_vector(9 downto 0);
    signal mulr_4_369 : std_logic_vector(9 downto 0);
    signal mulr_1_370 : std_logic_vector(9 downto 0);
    signal mulr_2_370 : std_logic_vector(9 downto 0);
    signal mulr_3_370 : std_logic_vector(9 downto 0);
    signal mulr_4_370 : std_logic_vector(9 downto 0);
    signal mulr_1_371 : std_logic_vector(9 downto 0);
    signal mulr_2_371 : std_logic_vector(9 downto 0);
    signal mulr_3_371 : std_logic_vector(9 downto 0);
    signal mulr_4_371 : std_logic_vector(9 downto 0);
    signal mulr_1_372 : std_logic_vector(9 downto 0);
    signal mulr_2_372 : std_logic_vector(9 downto 0);
    signal mulr_3_372 : std_logic_vector(9 downto 0);
    signal mulr_4_372 : std_logic_vector(9 downto 0);
    signal mulr_1_373 : std_logic_vector(9 downto 0);
    signal mulr_2_373 : std_logic_vector(9 downto 0);
    signal mulr_3_373 : std_logic_vector(9 downto 0);
    signal mulr_4_373 : std_logic_vector(9 downto 0);
    signal mulr_1_374 : std_logic_vector(9 downto 0);
    signal mulr_2_374 : std_logic_vector(9 downto 0);
    signal mulr_3_374 : std_logic_vector(9 downto 0);
    signal mulr_4_374 : std_logic_vector(9 downto 0);
    signal mulr_1_375 : std_logic_vector(9 downto 0);
    signal mulr_2_375 : std_logic_vector(9 downto 0);
    signal mulr_3_375 : std_logic_vector(9 downto 0);
    signal mulr_4_375 : std_logic_vector(9 downto 0);
    signal mulr_1_376 : std_logic_vector(9 downto 0);
    signal mulr_2_376 : std_logic_vector(9 downto 0);
    signal mulr_3_376 : std_logic_vector(9 downto 0);
    signal mulr_4_376 : std_logic_vector(9 downto 0);
    signal mulr_1_377 : std_logic_vector(9 downto 0);
    signal mulr_2_377 : std_logic_vector(9 downto 0);
    signal mulr_3_377 : std_logic_vector(9 downto 0);
    signal mulr_4_377 : std_logic_vector(9 downto 0);
    signal mulr_1_378 : std_logic_vector(9 downto 0);
    signal mulr_2_378 : std_logic_vector(9 downto 0);
    signal mulr_3_378 : std_logic_vector(9 downto 0);
    signal mulr_4_378 : std_logic_vector(9 downto 0);
    signal mulr_1_379 : std_logic_vector(9 downto 0);
    signal mulr_2_379 : std_logic_vector(9 downto 0);
    signal mulr_3_379 : std_logic_vector(9 downto 0);
    signal mulr_4_379 : std_logic_vector(9 downto 0);
    signal mulr_1_380 : std_logic_vector(9 downto 0);
    signal mulr_2_380 : std_logic_vector(9 downto 0);
    signal mulr_3_380 : std_logic_vector(9 downto 0);
    signal mulr_4_380 : std_logic_vector(9 downto 0);
    signal mulr_1_381 : std_logic_vector(9 downto 0);
    signal mulr_2_381 : std_logic_vector(9 downto 0);
    signal mulr_3_381 : std_logic_vector(9 downto 0);
    signal mulr_4_381 : std_logic_vector(9 downto 0);
    signal mulr_1_382 : std_logic_vector(9 downto 0);
    signal mulr_2_382 : std_logic_vector(9 downto 0);
    signal mulr_3_382 : std_logic_vector(9 downto 0);
    signal mulr_4_382 : std_logic_vector(9 downto 0);
    signal mulr_1_383 : std_logic_vector(9 downto 0);
    signal mulr_2_383 : std_logic_vector(9 downto 0);
    signal mulr_3_383 : std_logic_vector(9 downto 0);
    signal mulr_4_383 : std_logic_vector(9 downto 0);
    signal mulr_1_384 : std_logic_vector(9 downto 0);
    signal mulr_2_384 : std_logic_vector(9 downto 0);
    signal mulr_3_384 : std_logic_vector(9 downto 0);
    signal mulr_4_384 : std_logic_vector(9 downto 0);
    signal mulr_1_385 : std_logic_vector(9 downto 0);
    signal mulr_2_385 : std_logic_vector(9 downto 0);
    signal mulr_3_385 : std_logic_vector(9 downto 0);
    signal mulr_4_385 : std_logic_vector(9 downto 0);
    signal mulr_1_386 : std_logic_vector(9 downto 0);
    signal mulr_2_386 : std_logic_vector(9 downto 0);
    signal mulr_3_386 : std_logic_vector(9 downto 0);
    signal mulr_4_386 : std_logic_vector(9 downto 0);
    signal mulr_1_387 : std_logic_vector(9 downto 0);
    signal mulr_2_387 : std_logic_vector(9 downto 0);
    signal mulr_3_387 : std_logic_vector(9 downto 0);
    signal mulr_4_387 : std_logic_vector(9 downto 0);
    signal mulr_1_388 : std_logic_vector(9 downto 0);
    signal mulr_2_388 : std_logic_vector(9 downto 0);
    signal mulr_3_388 : std_logic_vector(9 downto 0);
    signal mulr_4_388 : std_logic_vector(9 downto 0);
    signal mulr_1_389 : std_logic_vector(9 downto 0);
    signal mulr_2_389 : std_logic_vector(9 downto 0);
    signal mulr_3_389 : std_logic_vector(9 downto 0);
    signal mulr_4_389 : std_logic_vector(9 downto 0);
    signal mulr_1_390 : std_logic_vector(9 downto 0);
    signal mulr_2_390 : std_logic_vector(9 downto 0);
    signal mulr_3_390 : std_logic_vector(9 downto 0);
    signal mulr_4_390 : std_logic_vector(9 downto 0);
    signal mulr_1_391 : std_logic_vector(9 downto 0);
    signal mulr_2_391 : std_logic_vector(9 downto 0);
    signal mulr_3_391 : std_logic_vector(9 downto 0);
    signal mulr_4_391 : std_logic_vector(9 downto 0);
    signal mulr_1_392 : std_logic_vector(9 downto 0);
    signal mulr_2_392 : std_logic_vector(9 downto 0);
    signal mulr_3_392 : std_logic_vector(9 downto 0);
    signal mulr_4_392 : std_logic_vector(9 downto 0);
    signal mulr_1_393 : std_logic_vector(9 downto 0);
    signal mulr_2_393 : std_logic_vector(9 downto 0);
    signal mulr_3_393 : std_logic_vector(9 downto 0);
    signal mulr_4_393 : std_logic_vector(9 downto 0);
    signal mulr_1_394 : std_logic_vector(9 downto 0);
    signal mulr_2_394 : std_logic_vector(9 downto 0);
    signal mulr_3_394 : std_logic_vector(9 downto 0);
    signal mulr_4_394 : std_logic_vector(9 downto 0);
    signal mulr_1_395 : std_logic_vector(9 downto 0);
    signal mulr_2_395 : std_logic_vector(9 downto 0);
    signal mulr_3_395 : std_logic_vector(9 downto 0);
    signal mulr_4_395 : std_logic_vector(9 downto 0);
    signal mulr_1_396 : std_logic_vector(9 downto 0);
    signal mulr_2_396 : std_logic_vector(9 downto 0);
    signal mulr_3_396 : std_logic_vector(9 downto 0);
    signal mulr_4_396 : std_logic_vector(9 downto 0);
    signal mulr_1_397 : std_logic_vector(9 downto 0);
    signal mulr_2_397 : std_logic_vector(9 downto 0);
    signal mulr_3_397 : std_logic_vector(9 downto 0);
    signal mulr_4_397 : std_logic_vector(9 downto 0);
    signal mulr_1_398 : std_logic_vector(9 downto 0);
    signal mulr_2_398 : std_logic_vector(9 downto 0);
    signal mulr_3_398 : std_logic_vector(9 downto 0);
    signal mulr_4_398 : std_logic_vector(9 downto 0);
    signal mulr_1_399 : std_logic_vector(9 downto 0);
    signal mulr_2_399 : std_logic_vector(9 downto 0);
    signal mulr_3_399 : std_logic_vector(9 downto 0);
    signal mulr_4_399 : std_logic_vector(9 downto 0);
    signal mulr_1_400 : std_logic_vector(9 downto 0);
    signal mulr_2_400 : std_logic_vector(9 downto 0);
    signal mulr_3_400 : std_logic_vector(9 downto 0);
    signal mulr_4_400 : std_logic_vector(9 downto 0);
    signal mulr_1_401 : std_logic_vector(9 downto 0);
    signal mulr_2_401 : std_logic_vector(9 downto 0);
    signal mulr_3_401 : std_logic_vector(9 downto 0);
    signal mulr_4_401 : std_logic_vector(9 downto 0);
    signal mulr_1_402 : std_logic_vector(9 downto 0);
    signal mulr_2_402 : std_logic_vector(9 downto 0);
    signal mulr_3_402 : std_logic_vector(9 downto 0);
    signal mulr_4_402 : std_logic_vector(9 downto 0);
    signal mulr_1_403 : std_logic_vector(9 downto 0);
    signal mulr_2_403 : std_logic_vector(9 downto 0);
    signal mulr_3_403 : std_logic_vector(9 downto 0);
    signal mulr_4_403 : std_logic_vector(9 downto 0);
    signal mulr_1_404 : std_logic_vector(9 downto 0);
    signal mulr_2_404 : std_logic_vector(9 downto 0);
    signal mulr_3_404 : std_logic_vector(9 downto 0);
    signal mulr_4_404 : std_logic_vector(9 downto 0);
    signal mulr_1_405 : std_logic_vector(9 downto 0);
    signal mulr_2_405 : std_logic_vector(9 downto 0);
    signal mulr_3_405 : std_logic_vector(9 downto 0);
    signal mulr_4_405 : std_logic_vector(9 downto 0);
    signal mulr_1_406 : std_logic_vector(9 downto 0);
    signal mulr_2_406 : std_logic_vector(9 downto 0);
    signal mulr_3_406 : std_logic_vector(9 downto 0);
    signal mulr_4_406 : std_logic_vector(9 downto 0);
    signal mulr_1_407 : std_logic_vector(9 downto 0);
    signal mulr_2_407 : std_logic_vector(9 downto 0);
    signal mulr_3_407 : std_logic_vector(9 downto 0);
    signal mulr_4_407 : std_logic_vector(9 downto 0);
    signal mulr_1_408 : std_logic_vector(9 downto 0);
    signal mulr_2_408 : std_logic_vector(9 downto 0);
    signal mulr_3_408 : std_logic_vector(9 downto 0);
    signal mulr_4_408 : std_logic_vector(9 downto 0);
    signal mulr_1_409 : std_logic_vector(9 downto 0);
    signal mulr_2_409 : std_logic_vector(9 downto 0);
    signal mulr_3_409 : std_logic_vector(9 downto 0);
    signal mulr_4_409 : std_logic_vector(9 downto 0);
    signal mulr_1_410 : std_logic_vector(9 downto 0);
    signal mulr_2_410 : std_logic_vector(9 downto 0);
    signal mulr_3_410 : std_logic_vector(9 downto 0);
    signal mulr_4_410 : std_logic_vector(9 downto 0);
    signal mulr_1_411 : std_logic_vector(9 downto 0);
    signal mulr_2_411 : std_logic_vector(9 downto 0);
    signal mulr_3_411 : std_logic_vector(9 downto 0);
    signal mulr_4_411 : std_logic_vector(9 downto 0);
    signal mulr_1_412 : std_logic_vector(9 downto 0);
    signal mulr_2_412 : std_logic_vector(9 downto 0);
    signal mulr_3_412 : std_logic_vector(9 downto 0);
    signal mulr_4_412 : std_logic_vector(9 downto 0);
    signal mulr_1_413 : std_logic_vector(9 downto 0);
    signal mulr_2_413 : std_logic_vector(9 downto 0);
    signal mulr_3_413 : std_logic_vector(9 downto 0);
    signal mulr_4_413 : std_logic_vector(9 downto 0);
    signal mulr_1_414 : std_logic_vector(9 downto 0);
    signal mulr_2_414 : std_logic_vector(9 downto 0);
    signal mulr_3_414 : std_logic_vector(9 downto 0);
    signal mulr_4_414 : std_logic_vector(9 downto 0);
    signal mulr_1_415 : std_logic_vector(9 downto 0);
    signal mulr_2_415 : std_logic_vector(9 downto 0);
    signal mulr_3_415 : std_logic_vector(9 downto 0);
    signal mulr_4_415 : std_logic_vector(9 downto 0);
    signal mulr_1_416 : std_logic_vector(9 downto 0);
    signal mulr_2_416 : std_logic_vector(9 downto 0);
    signal mulr_3_416 : std_logic_vector(9 downto 0);
    signal mulr_4_416 : std_logic_vector(9 downto 0);
    signal mulr_1_417 : std_logic_vector(9 downto 0);
    signal mulr_2_417 : std_logic_vector(9 downto 0);
    signal mulr_3_417 : std_logic_vector(9 downto 0);
    signal mulr_4_417 : std_logic_vector(9 downto 0);
    signal mulr_1_418 : std_logic_vector(9 downto 0);
    signal mulr_2_418 : std_logic_vector(9 downto 0);
    signal mulr_3_418 : std_logic_vector(9 downto 0);
    signal mulr_4_418 : std_logic_vector(9 downto 0);
    signal mulr_1_419 : std_logic_vector(9 downto 0);
    signal mulr_2_419 : std_logic_vector(9 downto 0);
    signal mulr_3_419 : std_logic_vector(9 downto 0);
    signal mulr_4_419 : std_logic_vector(9 downto 0);
    signal mulr_1_420 : std_logic_vector(9 downto 0);
    signal mulr_2_420 : std_logic_vector(9 downto 0);
    signal mulr_3_420 : std_logic_vector(9 downto 0);
    signal mulr_4_420 : std_logic_vector(9 downto 0);
    signal mulr_1_421 : std_logic_vector(9 downto 0);
    signal mulr_2_421 : std_logic_vector(9 downto 0);
    signal mulr_3_421 : std_logic_vector(9 downto 0);
    signal mulr_4_421 : std_logic_vector(9 downto 0);
    signal mulr_1_422 : std_logic_vector(9 downto 0);
    signal mulr_2_422 : std_logic_vector(9 downto 0);
    signal mulr_3_422 : std_logic_vector(9 downto 0);
    signal mulr_4_422 : std_logic_vector(9 downto 0);
    signal mulr_1_423 : std_logic_vector(9 downto 0);
    signal mulr_2_423 : std_logic_vector(9 downto 0);
    signal mulr_3_423 : std_logic_vector(9 downto 0);
    signal mulr_4_423 : std_logic_vector(9 downto 0);
    signal mulr_1_424 : std_logic_vector(9 downto 0);
    signal mulr_2_424 : std_logic_vector(9 downto 0);
    signal mulr_3_424 : std_logic_vector(9 downto 0);
    signal mulr_4_424 : std_logic_vector(9 downto 0);
    signal mulr_1_425 : std_logic_vector(9 downto 0);
    signal mulr_2_425 : std_logic_vector(9 downto 0);
    signal mulr_3_425 : std_logic_vector(9 downto 0);
    signal mulr_4_425 : std_logic_vector(9 downto 0);
    signal mulr_1_426 : std_logic_vector(9 downto 0);
    signal mulr_2_426 : std_logic_vector(9 downto 0);
    signal mulr_3_426 : std_logic_vector(9 downto 0);
    signal mulr_4_426 : std_logic_vector(9 downto 0);
    signal mulr_1_427 : std_logic_vector(9 downto 0);
    signal mulr_2_427 : std_logic_vector(9 downto 0);
    signal mulr_3_427 : std_logic_vector(9 downto 0);
    signal mulr_4_427 : std_logic_vector(9 downto 0);
    signal mulr_1_428 : std_logic_vector(9 downto 0);
    signal mulr_2_428 : std_logic_vector(9 downto 0);
    signal mulr_3_428 : std_logic_vector(9 downto 0);
    signal mulr_4_428 : std_logic_vector(9 downto 0);
    signal mulr_1_429 : std_logic_vector(9 downto 0);
    signal mulr_2_429 : std_logic_vector(9 downto 0);
    signal mulr_3_429 : std_logic_vector(9 downto 0);
    signal mulr_4_429 : std_logic_vector(9 downto 0);
    signal mulr_1_430 : std_logic_vector(9 downto 0);
    signal mulr_2_430 : std_logic_vector(9 downto 0);
    signal mulr_3_430 : std_logic_vector(9 downto 0);
    signal mulr_4_430 : std_logic_vector(9 downto 0);
    signal mulr_1_431 : std_logic_vector(9 downto 0);
    signal mulr_2_431 : std_logic_vector(9 downto 0);
    signal mulr_3_431 : std_logic_vector(9 downto 0);
    signal mulr_4_431 : std_logic_vector(9 downto 0);
    signal mulr_1_432 : std_logic_vector(9 downto 0);
    signal mulr_2_432 : std_logic_vector(9 downto 0);
    signal mulr_3_432 : std_logic_vector(9 downto 0);
    signal mulr_4_432 : std_logic_vector(9 downto 0);
    signal mulr_1_433 : std_logic_vector(9 downto 0);
    signal mulr_2_433 : std_logic_vector(9 downto 0);
    signal mulr_3_433 : std_logic_vector(9 downto 0);
    signal mulr_4_433 : std_logic_vector(9 downto 0);
    signal mulr_1_434 : std_logic_vector(9 downto 0);
    signal mulr_2_434 : std_logic_vector(9 downto 0);
    signal mulr_3_434 : std_logic_vector(9 downto 0);
    signal mulr_4_434 : std_logic_vector(9 downto 0);
    signal mulr_1_435 : std_logic_vector(9 downto 0);
    signal mulr_2_435 : std_logic_vector(9 downto 0);
    signal mulr_3_435 : std_logic_vector(9 downto 0);
    signal mulr_4_435 : std_logic_vector(9 downto 0);
    signal mulr_1_436 : std_logic_vector(9 downto 0);
    signal mulr_2_436 : std_logic_vector(9 downto 0);
    signal mulr_3_436 : std_logic_vector(9 downto 0);
    signal mulr_4_436 : std_logic_vector(9 downto 0);
    signal mulr_1_437 : std_logic_vector(9 downto 0);
    signal mulr_2_437 : std_logic_vector(9 downto 0);
    signal mulr_3_437 : std_logic_vector(9 downto 0);
    signal mulr_4_437 : std_logic_vector(9 downto 0);
    signal mulr_1_438 : std_logic_vector(9 downto 0);
    signal mulr_2_438 : std_logic_vector(9 downto 0);
    signal mulr_3_438 : std_logic_vector(9 downto 0);
    signal mulr_4_438 : std_logic_vector(9 downto 0);
    signal mulr_1_439 : std_logic_vector(9 downto 0);
    signal mulr_2_439 : std_logic_vector(9 downto 0);
    signal mulr_3_439 : std_logic_vector(9 downto 0);
    signal mulr_4_439 : std_logic_vector(9 downto 0);
    signal mulr_1_440 : std_logic_vector(9 downto 0);
    signal mulr_2_440 : std_logic_vector(9 downto 0);
    signal mulr_3_440 : std_logic_vector(9 downto 0);
    signal mulr_4_440 : std_logic_vector(9 downto 0);
    signal mulr_1_441 : std_logic_vector(9 downto 0);
    signal mulr_2_441 : std_logic_vector(9 downto 0);
    signal mulr_3_441 : std_logic_vector(9 downto 0);
    signal mulr_4_441 : std_logic_vector(9 downto 0);
    signal mulr_1_442 : std_logic_vector(9 downto 0);
    signal mulr_2_442 : std_logic_vector(9 downto 0);
    signal mulr_3_442 : std_logic_vector(9 downto 0);
    signal mulr_4_442 : std_logic_vector(9 downto 0);
    signal mulr_1_443 : std_logic_vector(9 downto 0);
    signal mulr_2_443 : std_logic_vector(9 downto 0);
    signal mulr_3_443 : std_logic_vector(9 downto 0);
    signal mulr_4_443 : std_logic_vector(9 downto 0);
    signal mulr_1_444 : std_logic_vector(9 downto 0);
    signal mulr_2_444 : std_logic_vector(9 downto 0);
    signal mulr_3_444 : std_logic_vector(9 downto 0);
    signal mulr_4_444 : std_logic_vector(9 downto 0);
    signal mulr_1_445 : std_logic_vector(9 downto 0);
    signal mulr_2_445 : std_logic_vector(9 downto 0);
    signal mulr_3_445 : std_logic_vector(9 downto 0);
    signal mulr_4_445 : std_logic_vector(9 downto 0);
    signal mulr_1_446 : std_logic_vector(9 downto 0);
    signal mulr_2_446 : std_logic_vector(9 downto 0);
    signal mulr_3_446 : std_logic_vector(9 downto 0);
    signal mulr_4_446 : std_logic_vector(9 downto 0);
    signal mulr_1_447 : std_logic_vector(9 downto 0);
    signal mulr_2_447 : std_logic_vector(9 downto 0);
    signal mulr_3_447 : std_logic_vector(9 downto 0);
    signal mulr_4_447 : std_logic_vector(9 downto 0);
    signal mulr_1_448 : std_logic_vector(9 downto 0);
    signal mulr_2_448 : std_logic_vector(9 downto 0);
    signal mulr_3_448 : std_logic_vector(9 downto 0);
    signal mulr_4_448 : std_logic_vector(9 downto 0);
    signal mulr_1_449 : std_logic_vector(9 downto 0);
    signal mulr_2_449 : std_logic_vector(9 downto 0);
    signal mulr_3_449 : std_logic_vector(9 downto 0);
    signal mulr_4_449 : std_logic_vector(9 downto 0);
    signal mulr_1_450 : std_logic_vector(9 downto 0);
    signal mulr_2_450 : std_logic_vector(9 downto 0);
    signal mulr_3_450 : std_logic_vector(9 downto 0);
    signal mulr_4_450 : std_logic_vector(9 downto 0);
    signal mulr_1_451 : std_logic_vector(9 downto 0);
    signal mulr_2_451 : std_logic_vector(9 downto 0);
    signal mulr_3_451 : std_logic_vector(9 downto 0);
    signal mulr_4_451 : std_logic_vector(9 downto 0);
    signal mulr_1_452 : std_logic_vector(9 downto 0);
    signal mulr_2_452 : std_logic_vector(9 downto 0);
    signal mulr_3_452 : std_logic_vector(9 downto 0);
    signal mulr_4_452 : std_logic_vector(9 downto 0);
    signal mulr_1_453 : std_logic_vector(9 downto 0);
    signal mulr_2_453 : std_logic_vector(9 downto 0);
    signal mulr_3_453 : std_logic_vector(9 downto 0);
    signal mulr_4_453 : std_logic_vector(9 downto 0);
    signal mulr_1_454 : std_logic_vector(9 downto 0);
    signal mulr_2_454 : std_logic_vector(9 downto 0);
    signal mulr_3_454 : std_logic_vector(9 downto 0);
    signal mulr_4_454 : std_logic_vector(9 downto 0);
    signal mulr_1_455 : std_logic_vector(9 downto 0);
    signal mulr_2_455 : std_logic_vector(9 downto 0);
    signal mulr_3_455 : std_logic_vector(9 downto 0);
    signal mulr_4_455 : std_logic_vector(9 downto 0);
    signal mulr_1_456 : std_logic_vector(9 downto 0);
    signal mulr_2_456 : std_logic_vector(9 downto 0);
    signal mulr_3_456 : std_logic_vector(9 downto 0);
    signal mulr_4_456 : std_logic_vector(9 downto 0);
    signal mulr_1_457 : std_logic_vector(9 downto 0);
    signal mulr_2_457 : std_logic_vector(9 downto 0);
    signal mulr_3_457 : std_logic_vector(9 downto 0);
    signal mulr_4_457 : std_logic_vector(9 downto 0);
    signal mulr_1_458 : std_logic_vector(9 downto 0);
    signal mulr_2_458 : std_logic_vector(9 downto 0);
    signal mulr_3_458 : std_logic_vector(9 downto 0);
    signal mulr_4_458 : std_logic_vector(9 downto 0);
    signal mulr_1_459 : std_logic_vector(9 downto 0);
    signal mulr_2_459 : std_logic_vector(9 downto 0);
    signal mulr_3_459 : std_logic_vector(9 downto 0);
    signal mulr_4_459 : std_logic_vector(9 downto 0);
    signal mulr_1_460 : std_logic_vector(9 downto 0);
    signal mulr_2_460 : std_logic_vector(9 downto 0);
    signal mulr_3_460 : std_logic_vector(9 downto 0);
    signal mulr_4_460 : std_logic_vector(9 downto 0);
    signal mulr_1_461 : std_logic_vector(9 downto 0);
    signal mulr_2_461 : std_logic_vector(9 downto 0);
    signal mulr_3_461 : std_logic_vector(9 downto 0);
    signal mulr_4_461 : std_logic_vector(9 downto 0);
    signal mulr_1_462 : std_logic_vector(9 downto 0);
    signal mulr_2_462 : std_logic_vector(9 downto 0);
    signal mulr_3_462 : std_logic_vector(9 downto 0);
    signal mulr_4_462 : std_logic_vector(9 downto 0);
    signal mulr_1_463 : std_logic_vector(9 downto 0);
    signal mulr_2_463 : std_logic_vector(9 downto 0);
    signal mulr_3_463 : std_logic_vector(9 downto 0);
    signal mulr_4_463 : std_logic_vector(9 downto 0);
    signal mulr_1_464 : std_logic_vector(9 downto 0);
    signal mulr_2_464 : std_logic_vector(9 downto 0);
    signal mulr_3_464 : std_logic_vector(9 downto 0);
    signal mulr_4_464 : std_logic_vector(9 downto 0);
    signal mulr_1_465 : std_logic_vector(9 downto 0);
    signal mulr_2_465 : std_logic_vector(9 downto 0);
    signal mulr_3_465 : std_logic_vector(9 downto 0);
    signal mulr_4_465 : std_logic_vector(9 downto 0);
    signal mulr_1_466 : std_logic_vector(9 downto 0);
    signal mulr_2_466 : std_logic_vector(9 downto 0);
    signal mulr_3_466 : std_logic_vector(9 downto 0);
    signal mulr_4_466 : std_logic_vector(9 downto 0);
    signal mulr_1_467 : std_logic_vector(9 downto 0);
    signal mulr_2_467 : std_logic_vector(9 downto 0);
    signal mulr_3_467 : std_logic_vector(9 downto 0);
    signal mulr_4_467 : std_logic_vector(9 downto 0);
    signal mulr_1_468 : std_logic_vector(9 downto 0);
    signal mulr_2_468 : std_logic_vector(9 downto 0);
    signal mulr_3_468 : std_logic_vector(9 downto 0);
    signal mulr_4_468 : std_logic_vector(9 downto 0);
    signal mulr_1_469 : std_logic_vector(9 downto 0);
    signal mulr_2_469 : std_logic_vector(9 downto 0);
    signal mulr_3_469 : std_logic_vector(9 downto 0);
    signal mulr_4_469 : std_logic_vector(9 downto 0);
    signal mulr_1_470 : std_logic_vector(9 downto 0);
    signal mulr_2_470 : std_logic_vector(9 downto 0);
    signal mulr_3_470 : std_logic_vector(9 downto 0);
    signal mulr_4_470 : std_logic_vector(9 downto 0);
    signal mulr_1_471 : std_logic_vector(9 downto 0);
    signal mulr_2_471 : std_logic_vector(9 downto 0);
    signal mulr_3_471 : std_logic_vector(9 downto 0);
    signal mulr_4_471 : std_logic_vector(9 downto 0);
    signal mulr_1_472 : std_logic_vector(9 downto 0);
    signal mulr_2_472 : std_logic_vector(9 downto 0);
    signal mulr_3_472 : std_logic_vector(9 downto 0);
    signal mulr_4_472 : std_logic_vector(9 downto 0);
    signal mulr_1_473 : std_logic_vector(9 downto 0);
    signal mulr_2_473 : std_logic_vector(9 downto 0);
    signal mulr_3_473 : std_logic_vector(9 downto 0);
    signal mulr_4_473 : std_logic_vector(9 downto 0);
    signal mulr_1_474 : std_logic_vector(9 downto 0);
    signal mulr_2_474 : std_logic_vector(9 downto 0);
    signal mulr_3_474 : std_logic_vector(9 downto 0);
    signal mulr_4_474 : std_logic_vector(9 downto 0);
    signal mulr_1_475 : std_logic_vector(9 downto 0);
    signal mulr_2_475 : std_logic_vector(9 downto 0);
    signal mulr_3_475 : std_logic_vector(9 downto 0);
    signal mulr_4_475 : std_logic_vector(9 downto 0);
    signal mulr_1_476 : std_logic_vector(9 downto 0);
    signal mulr_2_476 : std_logic_vector(9 downto 0);
    signal mulr_3_476 : std_logic_vector(9 downto 0);
    signal mulr_4_476 : std_logic_vector(9 downto 0);
    signal mulr_1_477 : std_logic_vector(9 downto 0);
    signal mulr_2_477 : std_logic_vector(9 downto 0);
    signal mulr_3_477 : std_logic_vector(9 downto 0);
    signal mulr_4_477 : std_logic_vector(9 downto 0);
    signal mulr_1_478 : std_logic_vector(9 downto 0);
    signal mulr_2_478 : std_logic_vector(9 downto 0);
    signal mulr_3_478 : std_logic_vector(9 downto 0);
    signal mulr_4_478 : std_logic_vector(9 downto 0);
    signal mulr_1_479 : std_logic_vector(9 downto 0);
    signal mulr_2_479 : std_logic_vector(9 downto 0);
    signal mulr_3_479 : std_logic_vector(9 downto 0);
    signal mulr_4_479 : std_logic_vector(9 downto 0);
    signal mulr_1_480 : std_logic_vector(9 downto 0);
    signal mulr_2_480 : std_logic_vector(9 downto 0);
    signal mulr_3_480 : std_logic_vector(9 downto 0);
    signal mulr_4_480 : std_logic_vector(9 downto 0);
    signal mulr_1_481 : std_logic_vector(9 downto 0);
    signal mulr_2_481 : std_logic_vector(9 downto 0);
    signal mulr_3_481 : std_logic_vector(9 downto 0);
    signal mulr_4_481 : std_logic_vector(9 downto 0);
    signal mulr_1_482 : std_logic_vector(9 downto 0);
    signal mulr_2_482 : std_logic_vector(9 downto 0);
    signal mulr_3_482 : std_logic_vector(9 downto 0);
    signal mulr_4_482 : std_logic_vector(9 downto 0);
    signal mulr_1_483 : std_logic_vector(9 downto 0);
    signal mulr_2_483 : std_logic_vector(9 downto 0);
    signal mulr_3_483 : std_logic_vector(9 downto 0);
    signal mulr_4_483 : std_logic_vector(9 downto 0);
    signal mulr_1_484 : std_logic_vector(9 downto 0);
    signal mulr_2_484 : std_logic_vector(9 downto 0);
    signal mulr_3_484 : std_logic_vector(9 downto 0);
    signal mulr_4_484 : std_logic_vector(9 downto 0);
    signal mulr_1_485 : std_logic_vector(9 downto 0);
    signal mulr_2_485 : std_logic_vector(9 downto 0);
    signal mulr_3_485 : std_logic_vector(9 downto 0);
    signal mulr_4_485 : std_logic_vector(9 downto 0);
    signal mulr_1_486 : std_logic_vector(9 downto 0);
    signal mulr_2_486 : std_logic_vector(9 downto 0);
    signal mulr_3_486 : std_logic_vector(9 downto 0);
    signal mulr_4_486 : std_logic_vector(9 downto 0);
    signal mulr_1_487 : std_logic_vector(9 downto 0);
    signal mulr_2_487 : std_logic_vector(9 downto 0);
    signal mulr_3_487 : std_logic_vector(9 downto 0);
    signal mulr_4_487 : std_logic_vector(9 downto 0);
    signal mulr_1_488 : std_logic_vector(9 downto 0);
    signal mulr_2_488 : std_logic_vector(9 downto 0);
    signal mulr_3_488 : std_logic_vector(9 downto 0);
    signal mulr_4_488 : std_logic_vector(9 downto 0);
    signal mulr_1_489 : std_logic_vector(9 downto 0);
    signal mulr_2_489 : std_logic_vector(9 downto 0);
    signal mulr_3_489 : std_logic_vector(9 downto 0);
    signal mulr_4_489 : std_logic_vector(9 downto 0);
    signal mulr_1_490 : std_logic_vector(9 downto 0);
    signal mulr_2_490 : std_logic_vector(9 downto 0);
    signal mulr_3_490 : std_logic_vector(9 downto 0);
    signal mulr_4_490 : std_logic_vector(9 downto 0);
    signal mulr_1_491 : std_logic_vector(9 downto 0);
    signal mulr_2_491 : std_logic_vector(9 downto 0);
    signal mulr_3_491 : std_logic_vector(9 downto 0);
    signal mulr_4_491 : std_logic_vector(9 downto 0);
    signal mulr_1_492 : std_logic_vector(9 downto 0);
    signal mulr_2_492 : std_logic_vector(9 downto 0);
    signal mulr_3_492 : std_logic_vector(9 downto 0);
    signal mulr_4_492 : std_logic_vector(9 downto 0);
    signal mulr_1_493 : std_logic_vector(9 downto 0);
    signal mulr_2_493 : std_logic_vector(9 downto 0);
    signal mulr_3_493 : std_logic_vector(9 downto 0);
    signal mulr_4_493 : std_logic_vector(9 downto 0);
    signal mulr_1_494 : std_logic_vector(9 downto 0);
    signal mulr_2_494 : std_logic_vector(9 downto 0);
    signal mulr_3_494 : std_logic_vector(9 downto 0);
    signal mulr_4_494 : std_logic_vector(9 downto 0);
    signal mulr_1_495 : std_logic_vector(9 downto 0);
    signal mulr_2_495 : std_logic_vector(9 downto 0);
    signal mulr_3_495 : std_logic_vector(9 downto 0);
    signal mulr_4_495 : std_logic_vector(9 downto 0);
    signal mulr_1_496 : std_logic_vector(9 downto 0);
    signal mulr_2_496 : std_logic_vector(9 downto 0);
    signal mulr_3_496 : std_logic_vector(9 downto 0);
    signal mulr_4_496 : std_logic_vector(9 downto 0);
    signal mulr_1_497 : std_logic_vector(9 downto 0);
    signal mulr_2_497 : std_logic_vector(9 downto 0);
    signal mulr_3_497 : std_logic_vector(9 downto 0);
    signal mulr_4_497 : std_logic_vector(9 downto 0);
    signal mulr_1_498 : std_logic_vector(9 downto 0);
    signal mulr_2_498 : std_logic_vector(9 downto 0);
    signal mulr_3_498 : std_logic_vector(9 downto 0);
    signal mulr_4_498 : std_logic_vector(9 downto 0);
    signal mulr_1_499 : std_logic_vector(9 downto 0);
    signal mulr_2_499 : std_logic_vector(9 downto 0);
    signal mulr_3_499 : std_logic_vector(9 downto 0);
    signal mulr_4_499 : std_logic_vector(9 downto 0);
    signal mulr_1_500 : std_logic_vector(9 downto 0);
    signal mulr_2_500 : std_logic_vector(9 downto 0);
    signal mulr_3_500 : std_logic_vector(9 downto 0);
    signal mulr_4_500 : std_logic_vector(9 downto 0);
    signal mulr_1_501 : std_logic_vector(9 downto 0);
    signal mulr_2_501 : std_logic_vector(9 downto 0);
    signal mulr_3_501 : std_logic_vector(9 downto 0);
    signal mulr_4_501 : std_logic_vector(9 downto 0);
    signal mulr_1_502 : std_logic_vector(9 downto 0);
    signal mulr_2_502 : std_logic_vector(9 downto 0);
    signal mulr_3_502 : std_logic_vector(9 downto 0);
    signal mulr_4_502 : std_logic_vector(9 downto 0);
    signal mulr_1_503 : std_logic_vector(9 downto 0);
    signal mulr_2_503 : std_logic_vector(9 downto 0);
    signal mulr_3_503 : std_logic_vector(9 downto 0);
    signal mulr_4_503 : std_logic_vector(9 downto 0);
    signal mulr_1_504 : std_logic_vector(9 downto 0);
    signal mulr_2_504 : std_logic_vector(9 downto 0);
    signal mulr_3_504 : std_logic_vector(9 downto 0);
    signal mulr_4_504 : std_logic_vector(9 downto 0);
    signal mulr_1_505 : std_logic_vector(9 downto 0);
    signal mulr_2_505 : std_logic_vector(9 downto 0);
    signal mulr_3_505 : std_logic_vector(9 downto 0);
    signal mulr_4_505 : std_logic_vector(9 downto 0);
    signal mulr_1_506 : std_logic_vector(9 downto 0);
    signal mulr_2_506 : std_logic_vector(9 downto 0);
    signal mulr_3_506 : std_logic_vector(9 downto 0);
    signal mulr_4_506 : std_logic_vector(9 downto 0);
    signal mulr_1_507 : std_logic_vector(9 downto 0);
    signal mulr_2_507 : std_logic_vector(9 downto 0);
    signal mulr_3_507 : std_logic_vector(9 downto 0);
    signal mulr_4_507 : std_logic_vector(9 downto 0);
    signal mulr_1_508 : std_logic_vector(9 downto 0);
    signal mulr_2_508 : std_logic_vector(9 downto 0);
    signal mulr_3_508 : std_logic_vector(9 downto 0);
    signal mulr_4_508 : std_logic_vector(9 downto 0);
    signal mulr_1_509 : std_logic_vector(9 downto 0);
    signal mulr_2_509 : std_logic_vector(9 downto 0);
    signal mulr_3_509 : std_logic_vector(9 downto 0);
    signal mulr_4_509 : std_logic_vector(9 downto 0);
    signal mulr_1_510 : std_logic_vector(9 downto 0);
    signal mulr_2_510 : std_logic_vector(9 downto 0);
    signal mulr_3_510 : std_logic_vector(9 downto 0);
    signal mulr_4_510 : std_logic_vector(9 downto 0);
    signal mulr_1_511 : std_logic_vector(9 downto 0);
    signal mulr_2_511 : std_logic_vector(9 downto 0);
    signal mulr_3_511 : std_logic_vector(9 downto 0);
    signal mulr_4_511 : std_logic_vector(9 downto 0);
    signal mulr_1_512 : std_logic_vector(9 downto 0);
    signal mulr_2_512 : std_logic_vector(9 downto 0);
    signal mulr_3_512 : std_logic_vector(9 downto 0);
    signal mulr_4_512 : std_logic_vector(9 downto 0);
    signal mulr_1_513 : std_logic_vector(9 downto 0);
    signal mulr_2_513 : std_logic_vector(9 downto 0);
    signal mulr_3_513 : std_logic_vector(9 downto 0);
    signal mulr_4_513 : std_logic_vector(9 downto 0);
    signal mulr_1_514 : std_logic_vector(9 downto 0);
    signal mulr_2_514 : std_logic_vector(9 downto 0);
    signal mulr_3_514 : std_logic_vector(9 downto 0);
    signal mulr_4_514 : std_logic_vector(9 downto 0);
    signal mulr_1_515 : std_logic_vector(9 downto 0);
    signal mulr_2_515 : std_logic_vector(9 downto 0);
    signal mulr_3_515 : std_logic_vector(9 downto 0);
    signal mulr_4_515 : std_logic_vector(9 downto 0);
    signal mulr_1_516 : std_logic_vector(9 downto 0);
    signal mulr_2_516 : std_logic_vector(9 downto 0);
    signal mulr_3_516 : std_logic_vector(9 downto 0);
    signal mulr_4_516 : std_logic_vector(9 downto 0);
    signal mulr_1_517 : std_logic_vector(9 downto 0);
    signal mulr_2_517 : std_logic_vector(9 downto 0);
    signal mulr_3_517 : std_logic_vector(9 downto 0);
    signal mulr_4_517 : std_logic_vector(9 downto 0);
    signal mulr_1_518 : std_logic_vector(9 downto 0);
    signal mulr_2_518 : std_logic_vector(9 downto 0);
    signal mulr_3_518 : std_logic_vector(9 downto 0);
    signal mulr_4_518 : std_logic_vector(9 downto 0);
    signal mulr_1_519 : std_logic_vector(9 downto 0);
    signal mulr_2_519 : std_logic_vector(9 downto 0);
    signal mulr_3_519 : std_logic_vector(9 downto 0);
    signal mulr_4_519 : std_logic_vector(9 downto 0);
    signal mulr_1_520 : std_logic_vector(9 downto 0);
    signal mulr_2_520 : std_logic_vector(9 downto 0);
    signal mulr_3_520 : std_logic_vector(9 downto 0);
    signal mulr_4_520 : std_logic_vector(9 downto 0);
    signal mulr_1_521 : std_logic_vector(9 downto 0);
    signal mulr_2_521 : std_logic_vector(9 downto 0);
    signal mulr_3_521 : std_logic_vector(9 downto 0);
    signal mulr_4_521 : std_logic_vector(9 downto 0);
    signal mulr_1_522 : std_logic_vector(9 downto 0);
    signal mulr_2_522 : std_logic_vector(9 downto 0);
    signal mulr_3_522 : std_logic_vector(9 downto 0);
    signal mulr_4_522 : std_logic_vector(9 downto 0);
    signal mulr_1_523 : std_logic_vector(9 downto 0);
    signal mulr_2_523 : std_logic_vector(9 downto 0);
    signal mulr_3_523 : std_logic_vector(9 downto 0);
    signal mulr_4_523 : std_logic_vector(9 downto 0);
    signal mulr_1_524 : std_logic_vector(9 downto 0);
    signal mulr_2_524 : std_logic_vector(9 downto 0);
    signal mulr_3_524 : std_logic_vector(9 downto 0);
    signal mulr_4_524 : std_logic_vector(9 downto 0);
    signal mulr_1_525 : std_logic_vector(9 downto 0);
    signal mulr_2_525 : std_logic_vector(9 downto 0);
    signal mulr_3_525 : std_logic_vector(9 downto 0);
    signal mulr_4_525 : std_logic_vector(9 downto 0);
    signal mulr_1_526 : std_logic_vector(9 downto 0);
    signal mulr_2_526 : std_logic_vector(9 downto 0);
    signal mulr_3_526 : std_logic_vector(9 downto 0);
    signal mulr_4_526 : std_logic_vector(9 downto 0);
    signal mulr_1_527 : std_logic_vector(9 downto 0);
    signal mulr_2_527 : std_logic_vector(9 downto 0);
    signal mulr_3_527 : std_logic_vector(9 downto 0);
    signal mulr_4_527 : std_logic_vector(9 downto 0);
    signal mulr_1_528 : std_logic_vector(9 downto 0);
    signal mulr_2_528 : std_logic_vector(9 downto 0);
    signal mulr_3_528 : std_logic_vector(9 downto 0);
    signal mulr_4_528 : std_logic_vector(9 downto 0);
    signal mulr_1_529 : std_logic_vector(9 downto 0);
    signal mulr_2_529 : std_logic_vector(9 downto 0);
    signal mulr_3_529 : std_logic_vector(9 downto 0);
    signal mulr_4_529 : std_logic_vector(9 downto 0);
    signal mulr_1_530 : std_logic_vector(9 downto 0);
    signal mulr_2_530 : std_logic_vector(9 downto 0);
    signal mulr_3_530 : std_logic_vector(9 downto 0);
    signal mulr_4_530 : std_logic_vector(9 downto 0);
    signal mulr_1_531 : std_logic_vector(9 downto 0);
    signal mulr_2_531 : std_logic_vector(9 downto 0);
    signal mulr_3_531 : std_logic_vector(9 downto 0);
    signal mulr_4_531 : std_logic_vector(9 downto 0);
    signal mulr_1_532 : std_logic_vector(9 downto 0);
    signal mulr_2_532 : std_logic_vector(9 downto 0);
    signal mulr_3_532 : std_logic_vector(9 downto 0);
    signal mulr_4_532 : std_logic_vector(9 downto 0);
    signal mulr_1_533 : std_logic_vector(9 downto 0);
    signal mulr_2_533 : std_logic_vector(9 downto 0);
    signal mulr_3_533 : std_logic_vector(9 downto 0);
    signal mulr_4_533 : std_logic_vector(9 downto 0);
    signal mulr_1_534 : std_logic_vector(9 downto 0);
    signal mulr_2_534 : std_logic_vector(9 downto 0);
    signal mulr_3_534 : std_logic_vector(9 downto 0);
    signal mulr_4_534 : std_logic_vector(9 downto 0);
    signal mulr_1_535 : std_logic_vector(9 downto 0);
    signal mulr_2_535 : std_logic_vector(9 downto 0);
    signal mulr_3_535 : std_logic_vector(9 downto 0);
    signal mulr_4_535 : std_logic_vector(9 downto 0);
    signal mulr_1_536 : std_logic_vector(9 downto 0);
    signal mulr_2_536 : std_logic_vector(9 downto 0);
    signal mulr_3_536 : std_logic_vector(9 downto 0);
    signal mulr_4_536 : std_logic_vector(9 downto 0);
    signal mulr_1_537 : std_logic_vector(9 downto 0);
    signal mulr_2_537 : std_logic_vector(9 downto 0);
    signal mulr_3_537 : std_logic_vector(9 downto 0);
    signal mulr_4_537 : std_logic_vector(9 downto 0);
    signal mulr_1_538 : std_logic_vector(9 downto 0);
    signal mulr_2_538 : std_logic_vector(9 downto 0);
    signal mulr_3_538 : std_logic_vector(9 downto 0);
    signal mulr_4_538 : std_logic_vector(9 downto 0);
    signal mulr_1_539 : std_logic_vector(9 downto 0);
    signal mulr_2_539 : std_logic_vector(9 downto 0);
    signal mulr_3_539 : std_logic_vector(9 downto 0);
    signal mulr_4_539 : std_logic_vector(9 downto 0);
    signal mulr_1_540 : std_logic_vector(9 downto 0);
    signal mulr_2_540 : std_logic_vector(9 downto 0);
    signal mulr_3_540 : std_logic_vector(9 downto 0);
    signal mulr_4_540 : std_logic_vector(9 downto 0);
    signal mulr_1_541 : std_logic_vector(9 downto 0);
    signal mulr_2_541 : std_logic_vector(9 downto 0);
    signal mulr_3_541 : std_logic_vector(9 downto 0);
    signal mulr_4_541 : std_logic_vector(9 downto 0);
    signal mulr_1_542 : std_logic_vector(9 downto 0);
    signal mulr_2_542 : std_logic_vector(9 downto 0);
    signal mulr_3_542 : std_logic_vector(9 downto 0);
    signal mulr_4_542 : std_logic_vector(9 downto 0);
    signal mulr_1_543 : std_logic_vector(9 downto 0);
    signal mulr_2_543 : std_logic_vector(9 downto 0);
    signal mulr_3_543 : std_logic_vector(9 downto 0);
    signal mulr_4_543 : std_logic_vector(9 downto 0);
    signal mulr_1_544 : std_logic_vector(9 downto 0);
    signal mulr_2_544 : std_logic_vector(9 downto 0);
    signal mulr_3_544 : std_logic_vector(9 downto 0);
    signal mulr_4_544 : std_logic_vector(9 downto 0);
    signal mulr_1_545 : std_logic_vector(9 downto 0);
    signal mulr_2_545 : std_logic_vector(9 downto 0);
    signal mulr_3_545 : std_logic_vector(9 downto 0);
    signal mulr_4_545 : std_logic_vector(9 downto 0);
    signal mulr_1_546 : std_logic_vector(9 downto 0);
    signal mulr_2_546 : std_logic_vector(9 downto 0);
    signal mulr_3_546 : std_logic_vector(9 downto 0);
    signal mulr_4_546 : std_logic_vector(9 downto 0);
    signal mulr_1_547 : std_logic_vector(9 downto 0);
    signal mulr_2_547 : std_logic_vector(9 downto 0);
    signal mulr_3_547 : std_logic_vector(9 downto 0);
    signal mulr_4_547 : std_logic_vector(9 downto 0);
    signal mulr_1_548 : std_logic_vector(9 downto 0);
    signal mulr_2_548 : std_logic_vector(9 downto 0);
    signal mulr_3_548 : std_logic_vector(9 downto 0);
    signal mulr_4_548 : std_logic_vector(9 downto 0);
    signal mulr_1_549 : std_logic_vector(9 downto 0);
    signal mulr_2_549 : std_logic_vector(9 downto 0);
    signal mulr_3_549 : std_logic_vector(9 downto 0);
    signal mulr_4_549 : std_logic_vector(9 downto 0);
    signal mulr_1_550 : std_logic_vector(9 downto 0);
    signal mulr_2_550 : std_logic_vector(9 downto 0);
    signal mulr_3_550 : std_logic_vector(9 downto 0);
    signal mulr_4_550 : std_logic_vector(9 downto 0);
    signal mulr_1_551 : std_logic_vector(9 downto 0);
    signal mulr_2_551 : std_logic_vector(9 downto 0);
    signal mulr_3_551 : std_logic_vector(9 downto 0);
    signal mulr_4_551 : std_logic_vector(9 downto 0);
    signal mulr_1_552 : std_logic_vector(9 downto 0);
    signal mulr_2_552 : std_logic_vector(9 downto 0);
    signal mulr_3_552 : std_logic_vector(9 downto 0);
    signal mulr_4_552 : std_logic_vector(9 downto 0);
    signal mulr_1_553 : std_logic_vector(9 downto 0);
    signal mulr_2_553 : std_logic_vector(9 downto 0);
    signal mulr_3_553 : std_logic_vector(9 downto 0);
    signal mulr_4_553 : std_logic_vector(9 downto 0);
    signal mulr_1_554 : std_logic_vector(9 downto 0);
    signal mulr_2_554 : std_logic_vector(9 downto 0);
    signal mulr_3_554 : std_logic_vector(9 downto 0);
    signal mulr_4_554 : std_logic_vector(9 downto 0);
    signal mulr_1_555 : std_logic_vector(9 downto 0);
    signal mulr_2_555 : std_logic_vector(9 downto 0);
    signal mulr_3_555 : std_logic_vector(9 downto 0);
    signal mulr_4_555 : std_logic_vector(9 downto 0);
    signal mulr_1_556 : std_logic_vector(9 downto 0);
    signal mulr_2_556 : std_logic_vector(9 downto 0);
    signal mulr_3_556 : std_logic_vector(9 downto 0);
    signal mulr_4_556 : std_logic_vector(9 downto 0);
    signal mulr_1_557 : std_logic_vector(9 downto 0);
    signal mulr_2_557 : std_logic_vector(9 downto 0);
    signal mulr_3_557 : std_logic_vector(9 downto 0);
    signal mulr_4_557 : std_logic_vector(9 downto 0);
    signal mulr_1_558 : std_logic_vector(9 downto 0);
    signal mulr_2_558 : std_logic_vector(9 downto 0);
    signal mulr_3_558 : std_logic_vector(9 downto 0);
    signal mulr_4_558 : std_logic_vector(9 downto 0);
    signal mulr_1_559 : std_logic_vector(9 downto 0);
    signal mulr_2_559 : std_logic_vector(9 downto 0);
    signal mulr_3_559 : std_logic_vector(9 downto 0);
    signal mulr_4_559 : std_logic_vector(9 downto 0);
    signal mulr_1_560 : std_logic_vector(9 downto 0);
    signal mulr_2_560 : std_logic_vector(9 downto 0);
    signal mulr_3_560 : std_logic_vector(9 downto 0);
    signal mulr_4_560 : std_logic_vector(9 downto 0);
    signal mulr_1_561 : std_logic_vector(9 downto 0);
    signal mulr_2_561 : std_logic_vector(9 downto 0);
    signal mulr_3_561 : std_logic_vector(9 downto 0);
    signal mulr_4_561 : std_logic_vector(9 downto 0);
    signal mulr_1_562 : std_logic_vector(9 downto 0);
    signal mulr_2_562 : std_logic_vector(9 downto 0);
    signal mulr_3_562 : std_logic_vector(9 downto 0);
    signal mulr_4_562 : std_logic_vector(9 downto 0);
    signal mulr_1_563 : std_logic_vector(9 downto 0);
    signal mulr_2_563 : std_logic_vector(9 downto 0);
    signal mulr_3_563 : std_logic_vector(9 downto 0);
    signal mulr_4_563 : std_logic_vector(9 downto 0);
    signal mulr_1_564 : std_logic_vector(9 downto 0);
    signal mulr_2_564 : std_logic_vector(9 downto 0);
    signal mulr_3_564 : std_logic_vector(9 downto 0);
    signal mulr_4_564 : std_logic_vector(9 downto 0);
    signal mulr_1_565 : std_logic_vector(9 downto 0);
    signal mulr_2_565 : std_logic_vector(9 downto 0);
    signal mulr_3_565 : std_logic_vector(9 downto 0);
    signal mulr_4_565 : std_logic_vector(9 downto 0);
    signal mulr_1_566 : std_logic_vector(9 downto 0);
    signal mulr_2_566 : std_logic_vector(9 downto 0);
    signal mulr_3_566 : std_logic_vector(9 downto 0);
    signal mulr_4_566 : std_logic_vector(9 downto 0);
    signal mulr_1_567 : std_logic_vector(9 downto 0);
    signal mulr_2_567 : std_logic_vector(9 downto 0);
    signal mulr_3_567 : std_logic_vector(9 downto 0);
    signal mulr_4_567 : std_logic_vector(9 downto 0);
    signal mulr_1_568 : std_logic_vector(9 downto 0);
    signal mulr_2_568 : std_logic_vector(9 downto 0);
    signal mulr_3_568 : std_logic_vector(9 downto 0);
    signal mulr_4_568 : std_logic_vector(9 downto 0);
    signal mulr_1_569 : std_logic_vector(9 downto 0);
    signal mulr_2_569 : std_logic_vector(9 downto 0);
    signal mulr_3_569 : std_logic_vector(9 downto 0);
    signal mulr_4_569 : std_logic_vector(9 downto 0);
    signal mulr_1_570 : std_logic_vector(9 downto 0);
    signal mulr_2_570 : std_logic_vector(9 downto 0);
    signal mulr_3_570 : std_logic_vector(9 downto 0);
    signal mulr_4_570 : std_logic_vector(9 downto 0);
    signal mulr_1_571 : std_logic_vector(9 downto 0);
    signal mulr_2_571 : std_logic_vector(9 downto 0);
    signal mulr_3_571 : std_logic_vector(9 downto 0);
    signal mulr_4_571 : std_logic_vector(9 downto 0);
    signal mulr_1_572 : std_logic_vector(9 downto 0);
    signal mulr_2_572 : std_logic_vector(9 downto 0);
    signal mulr_3_572 : std_logic_vector(9 downto 0);
    signal mulr_4_572 : std_logic_vector(9 downto 0);
    signal mulr_1_573 : std_logic_vector(9 downto 0);
    signal mulr_2_573 : std_logic_vector(9 downto 0);
    signal mulr_3_573 : std_logic_vector(9 downto 0);
    signal mulr_4_573 : std_logic_vector(9 downto 0);
    signal mulr_1_574 : std_logic_vector(9 downto 0);
    signal mulr_2_574 : std_logic_vector(9 downto 0);
    signal mulr_3_574 : std_logic_vector(9 downto 0);
    signal mulr_4_574 : std_logic_vector(9 downto 0);
    signal mulr_1_575 : std_logic_vector(9 downto 0);
    signal mulr_2_575 : std_logic_vector(9 downto 0);
    signal mulr_3_575 : std_logic_vector(9 downto 0);
    signal mulr_4_575 : std_logic_vector(9 downto 0);
    signal mulr_1_576 : std_logic_vector(9 downto 0);
    signal mulr_2_576 : std_logic_vector(9 downto 0);
    signal mulr_3_576 : std_logic_vector(9 downto 0);
    signal mulr_4_576 : std_logic_vector(9 downto 0);
    signal mulr_1_577 : std_logic_vector(9 downto 0);
    signal mulr_2_577 : std_logic_vector(9 downto 0);
    signal mulr_3_577 : std_logic_vector(9 downto 0);
    signal mulr_4_577 : std_logic_vector(9 downto 0);
    signal mulr_1_578 : std_logic_vector(9 downto 0);
    signal mulr_2_578 : std_logic_vector(9 downto 0);
    signal mulr_3_578 : std_logic_vector(9 downto 0);
    signal mulr_4_578 : std_logic_vector(9 downto 0);
    signal mulr_1_579 : std_logic_vector(9 downto 0);
    signal mulr_2_579 : std_logic_vector(9 downto 0);
    signal mulr_3_579 : std_logic_vector(9 downto 0);
    signal mulr_4_579 : std_logic_vector(9 downto 0);
    signal mulr_1_580 : std_logic_vector(9 downto 0);
    signal mulr_2_580 : std_logic_vector(9 downto 0);
    signal mulr_3_580 : std_logic_vector(9 downto 0);
    signal mulr_4_580 : std_logic_vector(9 downto 0);
    signal mulr_1_581 : std_logic_vector(9 downto 0);
    signal mulr_2_581 : std_logic_vector(9 downto 0);
    signal mulr_3_581 : std_logic_vector(9 downto 0);
    signal mulr_4_581 : std_logic_vector(9 downto 0);
    signal mulr_1_582 : std_logic_vector(9 downto 0);
    signal mulr_2_582 : std_logic_vector(9 downto 0);
    signal mulr_3_582 : std_logic_vector(9 downto 0);
    signal mulr_4_582 : std_logic_vector(9 downto 0);
    signal mulr_1_583 : std_logic_vector(9 downto 0);
    signal mulr_2_583 : std_logic_vector(9 downto 0);
    signal mulr_3_583 : std_logic_vector(9 downto 0);
    signal mulr_4_583 : std_logic_vector(9 downto 0);
    signal mulr_1_584 : std_logic_vector(9 downto 0);
    signal mulr_2_584 : std_logic_vector(9 downto 0);
    signal mulr_3_584 : std_logic_vector(9 downto 0);
    signal mulr_4_584 : std_logic_vector(9 downto 0);
    signal mulr_1_585 : std_logic_vector(9 downto 0);
    signal mulr_2_585 : std_logic_vector(9 downto 0);
    signal mulr_3_585 : std_logic_vector(9 downto 0);
    signal mulr_4_585 : std_logic_vector(9 downto 0);
    signal mulr_1_586 : std_logic_vector(9 downto 0);
    signal mulr_2_586 : std_logic_vector(9 downto 0);
    signal mulr_3_586 : std_logic_vector(9 downto 0);
    signal mulr_4_586 : std_logic_vector(9 downto 0);
    signal mulr_1_587 : std_logic_vector(9 downto 0);
    signal mulr_2_587 : std_logic_vector(9 downto 0);
    signal mulr_3_587 : std_logic_vector(9 downto 0);
    signal mulr_4_587 : std_logic_vector(9 downto 0);
    signal mulr_1_588 : std_logic_vector(9 downto 0);
    signal mulr_2_588 : std_logic_vector(9 downto 0);
    signal mulr_3_588 : std_logic_vector(9 downto 0);
    signal mulr_4_588 : std_logic_vector(9 downto 0);
    signal mulr_1_589 : std_logic_vector(9 downto 0);
    signal mulr_2_589 : std_logic_vector(9 downto 0);
    signal mulr_3_589 : std_logic_vector(9 downto 0);
    signal mulr_4_589 : std_logic_vector(9 downto 0);
    signal mulr_1_590 : std_logic_vector(9 downto 0);
    signal mulr_2_590 : std_logic_vector(9 downto 0);
    signal mulr_3_590 : std_logic_vector(9 downto 0);
    signal mulr_4_590 : std_logic_vector(9 downto 0);
    signal mulr_1_591 : std_logic_vector(9 downto 0);
    signal mulr_2_591 : std_logic_vector(9 downto 0);
    signal mulr_3_591 : std_logic_vector(9 downto 0);
    signal mulr_4_591 : std_logic_vector(9 downto 0);
    signal mulr_1_592 : std_logic_vector(9 downto 0);
    signal mulr_2_592 : std_logic_vector(9 downto 0);
    signal mulr_3_592 : std_logic_vector(9 downto 0);
    signal mulr_4_592 : std_logic_vector(9 downto 0);
    signal mulr_1_593 : std_logic_vector(9 downto 0);
    signal mulr_2_593 : std_logic_vector(9 downto 0);
    signal mulr_3_593 : std_logic_vector(9 downto 0);
    signal mulr_4_593 : std_logic_vector(9 downto 0);
    signal mulr_1_594 : std_logic_vector(9 downto 0);
    signal mulr_2_594 : std_logic_vector(9 downto 0);
    signal mulr_3_594 : std_logic_vector(9 downto 0);
    signal mulr_4_594 : std_logic_vector(9 downto 0);
    signal mulr_1_595 : std_logic_vector(9 downto 0);
    signal mulr_2_595 : std_logic_vector(9 downto 0);
    signal mulr_3_595 : std_logic_vector(9 downto 0);
    signal mulr_4_595 : std_logic_vector(9 downto 0);
    signal mulr_1_596 : std_logic_vector(9 downto 0);
    signal mulr_2_596 : std_logic_vector(9 downto 0);
    signal mulr_3_596 : std_logic_vector(9 downto 0);
    signal mulr_4_596 : std_logic_vector(9 downto 0);
    signal mulr_1_597 : std_logic_vector(9 downto 0);
    signal mulr_2_597 : std_logic_vector(9 downto 0);
    signal mulr_3_597 : std_logic_vector(9 downto 0);
    signal mulr_4_597 : std_logic_vector(9 downto 0);
    signal mulr_1_598 : std_logic_vector(9 downto 0);
    signal mulr_2_598 : std_logic_vector(9 downto 0);
    signal mulr_3_598 : std_logic_vector(9 downto 0);
    signal mulr_4_598 : std_logic_vector(9 downto 0);
    signal mulr_1_599 : std_logic_vector(9 downto 0);
    signal mulr_2_599 : std_logic_vector(9 downto 0);
    signal mulr_3_599 : std_logic_vector(9 downto 0);
    signal mulr_4_599 : std_logic_vector(9 downto 0);
    signal mulr_1_600 : std_logic_vector(9 downto 0);
    signal mulr_2_600 : std_logic_vector(9 downto 0);
    signal mulr_3_600 : std_logic_vector(9 downto 0);
    signal mulr_4_600 : std_logic_vector(9 downto 0);
    signal mulr_1_601 : std_logic_vector(9 downto 0);
    signal mulr_2_601 : std_logic_vector(9 downto 0);
    signal mulr_3_601 : std_logic_vector(9 downto 0);
    signal mulr_4_601 : std_logic_vector(9 downto 0);
    signal mulr_1_602 : std_logic_vector(9 downto 0);
    signal mulr_2_602 : std_logic_vector(9 downto 0);
    signal mulr_3_602 : std_logic_vector(9 downto 0);
    signal mulr_4_602 : std_logic_vector(9 downto 0);
    signal mulr_1_603 : std_logic_vector(9 downto 0);
    signal mulr_2_603 : std_logic_vector(9 downto 0);
    signal mulr_3_603 : std_logic_vector(9 downto 0);
    signal mulr_4_603 : std_logic_vector(9 downto 0);
    signal mulr_1_604 : std_logic_vector(9 downto 0);
    signal mulr_2_604 : std_logic_vector(9 downto 0);
    signal mulr_3_604 : std_logic_vector(9 downto 0);
    signal mulr_4_604 : std_logic_vector(9 downto 0);
    signal mulr_1_605 : std_logic_vector(9 downto 0);
    signal mulr_2_605 : std_logic_vector(9 downto 0);
    signal mulr_3_605 : std_logic_vector(9 downto 0);
    signal mulr_4_605 : std_logic_vector(9 downto 0);
    signal mulr_1_606 : std_logic_vector(9 downto 0);
    signal mulr_2_606 : std_logic_vector(9 downto 0);
    signal mulr_3_606 : std_logic_vector(9 downto 0);
    signal mulr_4_606 : std_logic_vector(9 downto 0);
    signal mulr_1_607 : std_logic_vector(9 downto 0);
    signal mulr_2_607 : std_logic_vector(9 downto 0);
    signal mulr_3_607 : std_logic_vector(9 downto 0);
    signal mulr_4_607 : std_logic_vector(9 downto 0);
    signal mulr_1_608 : std_logic_vector(9 downto 0);
    signal mulr_2_608 : std_logic_vector(9 downto 0);
    signal mulr_3_608 : std_logic_vector(9 downto 0);
    signal mulr_4_608 : std_logic_vector(9 downto 0);
    signal mulr_1_609 : std_logic_vector(9 downto 0);
    signal mulr_2_609 : std_logic_vector(9 downto 0);
    signal mulr_3_609 : std_logic_vector(9 downto 0);
    signal mulr_4_609 : std_logic_vector(9 downto 0);
    signal mulr_1_610 : std_logic_vector(9 downto 0);
    signal mulr_2_610 : std_logic_vector(9 downto 0);
    signal mulr_3_610 : std_logic_vector(9 downto 0);
    signal mulr_4_610 : std_logic_vector(9 downto 0);
    signal mulr_1_611 : std_logic_vector(9 downto 0);
    signal mulr_2_611 : std_logic_vector(9 downto 0);
    signal mulr_3_611 : std_logic_vector(9 downto 0);
    signal mulr_4_611 : std_logic_vector(9 downto 0);
    signal mulr_1_612 : std_logic_vector(9 downto 0);
    signal mulr_2_612 : std_logic_vector(9 downto 0);
    signal mulr_3_612 : std_logic_vector(9 downto 0);
    signal mulr_4_612 : std_logic_vector(9 downto 0);
    signal mulr_1_613 : std_logic_vector(9 downto 0);
    signal mulr_2_613 : std_logic_vector(9 downto 0);
    signal mulr_3_613 : std_logic_vector(9 downto 0);
    signal mulr_4_613 : std_logic_vector(9 downto 0);
    signal mulr_1_614 : std_logic_vector(9 downto 0);
    signal mulr_2_614 : std_logic_vector(9 downto 0);
    signal mulr_3_614 : std_logic_vector(9 downto 0);
    signal mulr_4_614 : std_logic_vector(9 downto 0);
    signal mulr_1_615 : std_logic_vector(9 downto 0);
    signal mulr_2_615 : std_logic_vector(9 downto 0);
    signal mulr_3_615 : std_logic_vector(9 downto 0);
    signal mulr_4_615 : std_logic_vector(9 downto 0);
    signal mulr_1_616 : std_logic_vector(9 downto 0);
    signal mulr_2_616 : std_logic_vector(9 downto 0);
    signal mulr_3_616 : std_logic_vector(9 downto 0);
    signal mulr_4_616 : std_logic_vector(9 downto 0);
    signal mulr_1_617 : std_logic_vector(9 downto 0);
    signal mulr_2_617 : std_logic_vector(9 downto 0);
    signal mulr_3_617 : std_logic_vector(9 downto 0);
    signal mulr_4_617 : std_logic_vector(9 downto 0);
    signal mulr_1_618 : std_logic_vector(9 downto 0);
    signal mulr_2_618 : std_logic_vector(9 downto 0);
    signal mulr_3_618 : std_logic_vector(9 downto 0);
    signal mulr_4_618 : std_logic_vector(9 downto 0);
    signal mulr_1_619 : std_logic_vector(9 downto 0);
    signal mulr_2_619 : std_logic_vector(9 downto 0);
    signal mulr_3_619 : std_logic_vector(9 downto 0);
    signal mulr_4_619 : std_logic_vector(9 downto 0);
    signal mulr_1_620 : std_logic_vector(9 downto 0);
    signal mulr_2_620 : std_logic_vector(9 downto 0);
    signal mulr_3_620 : std_logic_vector(9 downto 0);
    signal mulr_4_620 : std_logic_vector(9 downto 0);
    signal mulr_1_621 : std_logic_vector(9 downto 0);
    signal mulr_2_621 : std_logic_vector(9 downto 0);
    signal mulr_3_621 : std_logic_vector(9 downto 0);
    signal mulr_4_621 : std_logic_vector(9 downto 0);
    signal mulr_1_622 : std_logic_vector(9 downto 0);
    signal mulr_2_622 : std_logic_vector(9 downto 0);
    signal mulr_3_622 : std_logic_vector(9 downto 0);
    signal mulr_4_622 : std_logic_vector(9 downto 0);
    signal mulr_1_623 : std_logic_vector(9 downto 0);
    signal mulr_2_623 : std_logic_vector(9 downto 0);
    signal mulr_3_623 : std_logic_vector(9 downto 0);
    signal mulr_4_623 : std_logic_vector(9 downto 0);
    signal mulr_1_624 : std_logic_vector(9 downto 0);
    signal mulr_2_624 : std_logic_vector(9 downto 0);
    signal mulr_3_624 : std_logic_vector(9 downto 0);
    signal mulr_4_624 : std_logic_vector(9 downto 0);
    signal mulr_1_625 : std_logic_vector(9 downto 0);
    signal mulr_2_625 : std_logic_vector(9 downto 0);
    signal mulr_3_625 : std_logic_vector(9 downto 0);
    signal mulr_4_625 : std_logic_vector(9 downto 0);
    signal mulr_1_626 : std_logic_vector(9 downto 0);
    signal mulr_2_626 : std_logic_vector(9 downto 0);
    signal mulr_3_626 : std_logic_vector(9 downto 0);
    signal mulr_4_626 : std_logic_vector(9 downto 0);
    signal mulr_1_627 : std_logic_vector(9 downto 0);
    signal mulr_2_627 : std_logic_vector(9 downto 0);
    signal mulr_3_627 : std_logic_vector(9 downto 0);
    signal mulr_4_627 : std_logic_vector(9 downto 0);
    signal mulr_1_628 : std_logic_vector(9 downto 0);
    signal mulr_2_628 : std_logic_vector(9 downto 0);
    signal mulr_3_628 : std_logic_vector(9 downto 0);
    signal mulr_4_628 : std_logic_vector(9 downto 0);
    signal mulr_1_629 : std_logic_vector(9 downto 0);
    signal mulr_2_629 : std_logic_vector(9 downto 0);
    signal mulr_3_629 : std_logic_vector(9 downto 0);
    signal mulr_4_629 : std_logic_vector(9 downto 0);
    signal mulr_1_630 : std_logic_vector(9 downto 0);
    signal mulr_2_630 : std_logic_vector(9 downto 0);
    signal mulr_3_630 : std_logic_vector(9 downto 0);
    signal mulr_4_630 : std_logic_vector(9 downto 0);
    signal mulr_1_631 : std_logic_vector(9 downto 0);
    signal mulr_2_631 : std_logic_vector(9 downto 0);
    signal mulr_3_631 : std_logic_vector(9 downto 0);
    signal mulr_4_631 : std_logic_vector(9 downto 0);
    signal mulr_1_632 : std_logic_vector(9 downto 0);
    signal mulr_2_632 : std_logic_vector(9 downto 0);
    signal mulr_3_632 : std_logic_vector(9 downto 0);
    signal mulr_4_632 : std_logic_vector(9 downto 0);
    signal mulr_1_633 : std_logic_vector(9 downto 0);
    signal mulr_2_633 : std_logic_vector(9 downto 0);
    signal mulr_3_633 : std_logic_vector(9 downto 0);
    signal mulr_4_633 : std_logic_vector(9 downto 0);
    signal mulr_1_634 : std_logic_vector(9 downto 0);
    signal mulr_2_634 : std_logic_vector(9 downto 0);
    signal mulr_3_634 : std_logic_vector(9 downto 0);
    signal mulr_4_634 : std_logic_vector(9 downto 0);
    signal mulr_1_635 : std_logic_vector(9 downto 0);
    signal mulr_2_635 : std_logic_vector(9 downto 0);
    signal mulr_3_635 : std_logic_vector(9 downto 0);
    signal mulr_4_635 : std_logic_vector(9 downto 0);
    signal mulr_1_636 : std_logic_vector(9 downto 0);
    signal mulr_2_636 : std_logic_vector(9 downto 0);
    signal mulr_3_636 : std_logic_vector(9 downto 0);
    signal mulr_4_636 : std_logic_vector(9 downto 0);
    signal mulr_1_637 : std_logic_vector(9 downto 0);
    signal mulr_2_637 : std_logic_vector(9 downto 0);
    signal mulr_3_637 : std_logic_vector(9 downto 0);
    signal mulr_4_637 : std_logic_vector(9 downto 0);
    signal mulr_1_638 : std_logic_vector(9 downto 0);
    signal mulr_2_638 : std_logic_vector(9 downto 0);
    signal mulr_3_638 : std_logic_vector(9 downto 0);
    signal mulr_4_638 : std_logic_vector(9 downto 0);
    signal mulr_1_639 : std_logic_vector(9 downto 0);
    signal mulr_2_639 : std_logic_vector(9 downto 0);
    signal mulr_3_639 : std_logic_vector(9 downto 0);
    signal mulr_4_639 : std_logic_vector(9 downto 0);
    signal mulr_1_640 : std_logic_vector(9 downto 0);
    signal mulr_2_640 : std_logic_vector(9 downto 0);
    signal mulr_3_640 : std_logic_vector(9 downto 0);
    signal mulr_4_640 : std_logic_vector(9 downto 0);
    signal mulr_1_641 : std_logic_vector(9 downto 0);
    signal mulr_2_641 : std_logic_vector(9 downto 0);
    signal mulr_3_641 : std_logic_vector(9 downto 0);
    signal mulr_4_641 : std_logic_vector(9 downto 0);
    signal mulr_1_642 : std_logic_vector(9 downto 0);
    signal mulr_2_642 : std_logic_vector(9 downto 0);
    signal mulr_3_642 : std_logic_vector(9 downto 0);
    signal mulr_4_642 : std_logic_vector(9 downto 0);
    signal mulr_1_643 : std_logic_vector(9 downto 0);
    signal mulr_2_643 : std_logic_vector(9 downto 0);
    signal mulr_3_643 : std_logic_vector(9 downto 0);
    signal mulr_4_643 : std_logic_vector(9 downto 0);
    signal mulr_1_644 : std_logic_vector(9 downto 0);
    signal mulr_2_644 : std_logic_vector(9 downto 0);
    signal mulr_3_644 : std_logic_vector(9 downto 0);
    signal mulr_4_644 : std_logic_vector(9 downto 0);
    signal mulr_1_645 : std_logic_vector(9 downto 0);
    signal mulr_2_645 : std_logic_vector(9 downto 0);
    signal mulr_3_645 : std_logic_vector(9 downto 0);
    signal mulr_4_645 : std_logic_vector(9 downto 0);
    signal mulr_1_646 : std_logic_vector(9 downto 0);
    signal mulr_2_646 : std_logic_vector(9 downto 0);
    signal mulr_3_646 : std_logic_vector(9 downto 0);
    signal mulr_4_646 : std_logic_vector(9 downto 0);
    signal mulr_1_647 : std_logic_vector(9 downto 0);
    signal mulr_2_647 : std_logic_vector(9 downto 0);
    signal mulr_3_647 : std_logic_vector(9 downto 0);
    signal mulr_4_647 : std_logic_vector(9 downto 0);
    signal mulr_1_648 : std_logic_vector(9 downto 0);
    signal mulr_2_648 : std_logic_vector(9 downto 0);
    signal mulr_3_648 : std_logic_vector(9 downto 0);
    signal mulr_4_648 : std_logic_vector(9 downto 0);
    signal mulr_1_649 : std_logic_vector(9 downto 0);
    signal mulr_2_649 : std_logic_vector(9 downto 0);
    signal mulr_3_649 : std_logic_vector(9 downto 0);
    signal mulr_4_649 : std_logic_vector(9 downto 0);
    signal mulr_1_650 : std_logic_vector(9 downto 0);
    signal mulr_2_650 : std_logic_vector(9 downto 0);
    signal mulr_3_650 : std_logic_vector(9 downto 0);
    signal mulr_4_650 : std_logic_vector(9 downto 0);
    signal mulr_1_651 : std_logic_vector(9 downto 0);
    signal mulr_2_651 : std_logic_vector(9 downto 0);
    signal mulr_3_651 : std_logic_vector(9 downto 0);
    signal mulr_4_651 : std_logic_vector(9 downto 0);
    signal mulr_1_652 : std_logic_vector(9 downto 0);
    signal mulr_2_652 : std_logic_vector(9 downto 0);
    signal mulr_3_652 : std_logic_vector(9 downto 0);
    signal mulr_4_652 : std_logic_vector(9 downto 0);
    signal mulr_1_653 : std_logic_vector(9 downto 0);
    signal mulr_2_653 : std_logic_vector(9 downto 0);
    signal mulr_3_653 : std_logic_vector(9 downto 0);
    signal mulr_4_653 : std_logic_vector(9 downto 0);
    signal mulr_1_654 : std_logic_vector(9 downto 0);
    signal mulr_2_654 : std_logic_vector(9 downto 0);
    signal mulr_3_654 : std_logic_vector(9 downto 0);
    signal mulr_4_654 : std_logic_vector(9 downto 0);
    signal mulr_1_655 : std_logic_vector(9 downto 0);
    signal mulr_2_655 : std_logic_vector(9 downto 0);
    signal mulr_3_655 : std_logic_vector(9 downto 0);
    signal mulr_4_655 : std_logic_vector(9 downto 0);
    signal mulr_1_656 : std_logic_vector(9 downto 0);
    signal mulr_2_656 : std_logic_vector(9 downto 0);
    signal mulr_3_656 : std_logic_vector(9 downto 0);
    signal mulr_4_656 : std_logic_vector(9 downto 0);
    signal mulr_1_657 : std_logic_vector(9 downto 0);
    signal mulr_2_657 : std_logic_vector(9 downto 0);
    signal mulr_3_657 : std_logic_vector(9 downto 0);
    signal mulr_4_657 : std_logic_vector(9 downto 0);
    signal mulr_1_658 : std_logic_vector(9 downto 0);
    signal mulr_2_658 : std_logic_vector(9 downto 0);
    signal mulr_3_658 : std_logic_vector(9 downto 0);
    signal mulr_4_658 : std_logic_vector(9 downto 0);
    signal mulr_1_659 : std_logic_vector(9 downto 0);
    signal mulr_2_659 : std_logic_vector(9 downto 0);
    signal mulr_3_659 : std_logic_vector(9 downto 0);
    signal mulr_4_659 : std_logic_vector(9 downto 0);
    signal mulr_1_660 : std_logic_vector(9 downto 0);
    signal mulr_2_660 : std_logic_vector(9 downto 0);
    signal mulr_3_660 : std_logic_vector(9 downto 0);
    signal mulr_4_660 : std_logic_vector(9 downto 0);
    signal mulr_1_661 : std_logic_vector(9 downto 0);
    signal mulr_2_661 : std_logic_vector(9 downto 0);
    signal mulr_3_661 : std_logic_vector(9 downto 0);
    signal mulr_4_661 : std_logic_vector(9 downto 0);
    signal mulr_1_662 : std_logic_vector(9 downto 0);
    signal mulr_2_662 : std_logic_vector(9 downto 0);
    signal mulr_3_662 : std_logic_vector(9 downto 0);
    signal mulr_4_662 : std_logic_vector(9 downto 0);
    signal mulr_1_663 : std_logic_vector(9 downto 0);
    signal mulr_2_663 : std_logic_vector(9 downto 0);
    signal mulr_3_663 : std_logic_vector(9 downto 0);
    signal mulr_4_663 : std_logic_vector(9 downto 0);
    signal mulr_1_664 : std_logic_vector(9 downto 0);
    signal mulr_2_664 : std_logic_vector(9 downto 0);
    signal mulr_3_664 : std_logic_vector(9 downto 0);
    signal mulr_4_664 : std_logic_vector(9 downto 0);
    signal mulr_1_665 : std_logic_vector(9 downto 0);
    signal mulr_2_665 : std_logic_vector(9 downto 0);
    signal mulr_3_665 : std_logic_vector(9 downto 0);
    signal mulr_4_665 : std_logic_vector(9 downto 0);
    signal mulr_1_666 : std_logic_vector(9 downto 0);
    signal mulr_2_666 : std_logic_vector(9 downto 0);
    signal mulr_3_666 : std_logic_vector(9 downto 0);
    signal mulr_4_666 : std_logic_vector(9 downto 0);
    signal mulr_1_667 : std_logic_vector(9 downto 0);
    signal mulr_2_667 : std_logic_vector(9 downto 0);
    signal mulr_3_667 : std_logic_vector(9 downto 0);
    signal mulr_4_667 : std_logic_vector(9 downto 0);
    signal mulr_1_668 : std_logic_vector(9 downto 0);
    signal mulr_2_668 : std_logic_vector(9 downto 0);
    signal mulr_3_668 : std_logic_vector(9 downto 0);
    signal mulr_4_668 : std_logic_vector(9 downto 0);
    signal mulr_1_669 : std_logic_vector(9 downto 0);
    signal mulr_2_669 : std_logic_vector(9 downto 0);
    signal mulr_3_669 : std_logic_vector(9 downto 0);
    signal mulr_4_669 : std_logic_vector(9 downto 0);
    signal mulr_1_670 : std_logic_vector(9 downto 0);
    signal mulr_2_670 : std_logic_vector(9 downto 0);
    signal mulr_3_670 : std_logic_vector(9 downto 0);
    signal mulr_4_670 : std_logic_vector(9 downto 0);
    signal mulr_1_671 : std_logic_vector(9 downto 0);
    signal mulr_2_671 : std_logic_vector(9 downto 0);
    signal mulr_3_671 : std_logic_vector(9 downto 0);
    signal mulr_4_671 : std_logic_vector(9 downto 0);
    signal mulr_1_672 : std_logic_vector(9 downto 0);
    signal mulr_2_672 : std_logic_vector(9 downto 0);
    signal mulr_3_672 : std_logic_vector(9 downto 0);
    signal mulr_4_672 : std_logic_vector(9 downto 0);
    signal mulr_1_673 : std_logic_vector(9 downto 0);
    signal mulr_2_673 : std_logic_vector(9 downto 0);
    signal mulr_3_673 : std_logic_vector(9 downto 0);
    signal mulr_4_673 : std_logic_vector(9 downto 0);
    signal mulr_1_674 : std_logic_vector(9 downto 0);
    signal mulr_2_674 : std_logic_vector(9 downto 0);
    signal mulr_3_674 : std_logic_vector(9 downto 0);
    signal mulr_4_674 : std_logic_vector(9 downto 0);
    signal mulr_1_675 : std_logic_vector(9 downto 0);
    signal mulr_2_675 : std_logic_vector(9 downto 0);
    signal mulr_3_675 : std_logic_vector(9 downto 0);
    signal mulr_4_675 : std_logic_vector(9 downto 0);
    signal mulr_1_676 : std_logic_vector(9 downto 0);
    signal mulr_2_676 : std_logic_vector(9 downto 0);
    signal mulr_3_676 : std_logic_vector(9 downto 0);
    signal mulr_4_676 : std_logic_vector(9 downto 0);
    signal mulr_1_677 : std_logic_vector(9 downto 0);
    signal mulr_2_677 : std_logic_vector(9 downto 0);
    signal mulr_3_677 : std_logic_vector(9 downto 0);
    signal mulr_4_677 : std_logic_vector(9 downto 0);
    signal mulr_1_678 : std_logic_vector(9 downto 0);
    signal mulr_2_678 : std_logic_vector(9 downto 0);
    signal mulr_3_678 : std_logic_vector(9 downto 0);
    signal mulr_4_678 : std_logic_vector(9 downto 0);
    signal mulr_1_679 : std_logic_vector(9 downto 0);
    signal mulr_2_679 : std_logic_vector(9 downto 0);
    signal mulr_3_679 : std_logic_vector(9 downto 0);
    signal mulr_4_679 : std_logic_vector(9 downto 0);
    signal mulr_1_680 : std_logic_vector(9 downto 0);
    signal mulr_2_680 : std_logic_vector(9 downto 0);
    signal mulr_3_680 : std_logic_vector(9 downto 0);
    signal mulr_4_680 : std_logic_vector(9 downto 0);
    signal mulr_1_681 : std_logic_vector(9 downto 0);
    signal mulr_2_681 : std_logic_vector(9 downto 0);
    signal mulr_3_681 : std_logic_vector(9 downto 0);
    signal mulr_4_681 : std_logic_vector(9 downto 0);
    signal mulr_1_682 : std_logic_vector(9 downto 0);
    signal mulr_2_682 : std_logic_vector(9 downto 0);
    signal mulr_3_682 : std_logic_vector(9 downto 0);
    signal mulr_4_682 : std_logic_vector(9 downto 0);
    signal mulr_1_683 : std_logic_vector(9 downto 0);
    signal mulr_2_683 : std_logic_vector(9 downto 0);
    signal mulr_3_683 : std_logic_vector(9 downto 0);
    signal mulr_4_683 : std_logic_vector(9 downto 0);
    signal mulr_1_684 : std_logic_vector(9 downto 0);
    signal mulr_2_684 : std_logic_vector(9 downto 0);
    signal mulr_3_684 : std_logic_vector(9 downto 0);
    signal mulr_4_684 : std_logic_vector(9 downto 0);
    signal mulr_1_685 : std_logic_vector(9 downto 0);
    signal mulr_2_685 : std_logic_vector(9 downto 0);
    signal mulr_3_685 : std_logic_vector(9 downto 0);
    signal mulr_4_685 : std_logic_vector(9 downto 0);
    signal mulr_1_686 : std_logic_vector(9 downto 0);
    signal mulr_2_686 : std_logic_vector(9 downto 0);
    signal mulr_3_686 : std_logic_vector(9 downto 0);
    signal mulr_4_686 : std_logic_vector(9 downto 0);
    signal mulr_1_687 : std_logic_vector(9 downto 0);
    signal mulr_2_687 : std_logic_vector(9 downto 0);
    signal mulr_3_687 : std_logic_vector(9 downto 0);
    signal mulr_4_687 : std_logic_vector(9 downto 0);
    signal mulr_1_688 : std_logic_vector(9 downto 0);
    signal mulr_2_688 : std_logic_vector(9 downto 0);
    signal mulr_3_688 : std_logic_vector(9 downto 0);
    signal mulr_4_688 : std_logic_vector(9 downto 0);
    signal mulr_1_689 : std_logic_vector(9 downto 0);
    signal mulr_2_689 : std_logic_vector(9 downto 0);
    signal mulr_3_689 : std_logic_vector(9 downto 0);
    signal mulr_4_689 : std_logic_vector(9 downto 0);
    signal mulr_1_690 : std_logic_vector(9 downto 0);
    signal mulr_2_690 : std_logic_vector(9 downto 0);
    signal mulr_3_690 : std_logic_vector(9 downto 0);
    signal mulr_4_690 : std_logic_vector(9 downto 0);
    signal mulr_1_691 : std_logic_vector(9 downto 0);
    signal mulr_2_691 : std_logic_vector(9 downto 0);
    signal mulr_3_691 : std_logic_vector(9 downto 0);
    signal mulr_4_691 : std_logic_vector(9 downto 0);
    signal mulr_1_692 : std_logic_vector(9 downto 0);
    signal mulr_2_692 : std_logic_vector(9 downto 0);
    signal mulr_3_692 : std_logic_vector(9 downto 0);
    signal mulr_4_692 : std_logic_vector(9 downto 0);
    signal mulr_1_693 : std_logic_vector(9 downto 0);
    signal mulr_2_693 : std_logic_vector(9 downto 0);
    signal mulr_3_693 : std_logic_vector(9 downto 0);
    signal mulr_4_693 : std_logic_vector(9 downto 0);
    signal mulr_1_694 : std_logic_vector(9 downto 0);
    signal mulr_2_694 : std_logic_vector(9 downto 0);
    signal mulr_3_694 : std_logic_vector(9 downto 0);
    signal mulr_4_694 : std_logic_vector(9 downto 0);
    signal mulr_1_695 : std_logic_vector(9 downto 0);
    signal mulr_2_695 : std_logic_vector(9 downto 0);
    signal mulr_3_695 : std_logic_vector(9 downto 0);
    signal mulr_4_695 : std_logic_vector(9 downto 0);
    signal mulr_1_696 : std_logic_vector(9 downto 0);
    signal mulr_2_696 : std_logic_vector(9 downto 0);
    signal mulr_3_696 : std_logic_vector(9 downto 0);
    signal mulr_4_696 : std_logic_vector(9 downto 0);
    signal mulr_1_697 : std_logic_vector(9 downto 0);
    signal mulr_2_697 : std_logic_vector(9 downto 0);
    signal mulr_3_697 : std_logic_vector(9 downto 0);
    signal mulr_4_697 : std_logic_vector(9 downto 0);
    signal mulr_1_698 : std_logic_vector(9 downto 0);
    signal mulr_2_698 : std_logic_vector(9 downto 0);
    signal mulr_3_698 : std_logic_vector(9 downto 0);
    signal mulr_4_698 : std_logic_vector(9 downto 0);
    signal mulr_1_699 : std_logic_vector(9 downto 0);
    signal mulr_2_699 : std_logic_vector(9 downto 0);
    signal mulr_3_699 : std_logic_vector(9 downto 0);
    signal mulr_4_699 : std_logic_vector(9 downto 0);
    signal mulr_1_700 : std_logic_vector(9 downto 0);
    signal mulr_2_700 : std_logic_vector(9 downto 0);
    signal mulr_3_700 : std_logic_vector(9 downto 0);
    signal mulr_4_700 : std_logic_vector(9 downto 0);
    signal mulr_1_701 : std_logic_vector(9 downto 0);
    signal mulr_2_701 : std_logic_vector(9 downto 0);
    signal mulr_3_701 : std_logic_vector(9 downto 0);
    signal mulr_4_701 : std_logic_vector(9 downto 0);
    signal mulr_1_702 : std_logic_vector(9 downto 0);
    signal mulr_2_702 : std_logic_vector(9 downto 0);
    signal mulr_3_702 : std_logic_vector(9 downto 0);
    signal mulr_4_702 : std_logic_vector(9 downto 0);
    signal mulr_1_703 : std_logic_vector(9 downto 0);
    signal mulr_2_703 : std_logic_vector(9 downto 0);
    signal mulr_3_703 : std_logic_vector(9 downto 0);
    signal mulr_4_703 : std_logic_vector(9 downto 0);
    signal mulr_1_704 : std_logic_vector(9 downto 0);
    signal mulr_2_704 : std_logic_vector(9 downto 0);
    signal mulr_3_704 : std_logic_vector(9 downto 0);
    signal mulr_4_704 : std_logic_vector(9 downto 0);
    signal mulr_1_705 : std_logic_vector(9 downto 0);
    signal mulr_2_705 : std_logic_vector(9 downto 0);
    signal mulr_3_705 : std_logic_vector(9 downto 0);
    signal mulr_4_705 : std_logic_vector(9 downto 0);
    signal mulr_1_706 : std_logic_vector(9 downto 0);
    signal mulr_2_706 : std_logic_vector(9 downto 0);
    signal mulr_3_706 : std_logic_vector(9 downto 0);
    signal mulr_4_706 : std_logic_vector(9 downto 0);
    signal mulr_1_707 : std_logic_vector(9 downto 0);
    signal mulr_2_707 : std_logic_vector(9 downto 0);
    signal mulr_3_707 : std_logic_vector(9 downto 0);
    signal mulr_4_707 : std_logic_vector(9 downto 0);
    signal mulr_1_708 : std_logic_vector(9 downto 0);
    signal mulr_2_708 : std_logic_vector(9 downto 0);
    signal mulr_3_708 : std_logic_vector(9 downto 0);
    signal mulr_4_708 : std_logic_vector(9 downto 0);
    signal mulr_1_709 : std_logic_vector(9 downto 0);
    signal mulr_2_709 : std_logic_vector(9 downto 0);
    signal mulr_3_709 : std_logic_vector(9 downto 0);
    signal mulr_4_709 : std_logic_vector(9 downto 0);
    signal mulr_1_710 : std_logic_vector(9 downto 0);
    signal mulr_2_710 : std_logic_vector(9 downto 0);
    signal mulr_3_710 : std_logic_vector(9 downto 0);
    signal mulr_4_710 : std_logic_vector(9 downto 0);
    signal mulr_1_711 : std_logic_vector(9 downto 0);
    signal mulr_2_711 : std_logic_vector(9 downto 0);
    signal mulr_3_711 : std_logic_vector(9 downto 0);
    signal mulr_4_711 : std_logic_vector(9 downto 0);
    signal mulr_1_712 : std_logic_vector(9 downto 0);
    signal mulr_2_712 : std_logic_vector(9 downto 0);
    signal mulr_3_712 : std_logic_vector(9 downto 0);
    signal mulr_4_712 : std_logic_vector(9 downto 0);
    signal mulr_1_713 : std_logic_vector(9 downto 0);
    signal mulr_2_713 : std_logic_vector(9 downto 0);
    signal mulr_3_713 : std_logic_vector(9 downto 0);
    signal mulr_4_713 : std_logic_vector(9 downto 0);
    signal mulr_1_714 : std_logic_vector(9 downto 0);
    signal mulr_2_714 : std_logic_vector(9 downto 0);
    signal mulr_3_714 : std_logic_vector(9 downto 0);
    signal mulr_4_714 : std_logic_vector(9 downto 0);
    signal mulr_1_715 : std_logic_vector(9 downto 0);
    signal mulr_2_715 : std_logic_vector(9 downto 0);
    signal mulr_3_715 : std_logic_vector(9 downto 0);
    signal mulr_4_715 : std_logic_vector(9 downto 0);
    signal mulr_1_716 : std_logic_vector(9 downto 0);
    signal mulr_2_716 : std_logic_vector(9 downto 0);
    signal mulr_3_716 : std_logic_vector(9 downto 0);
    signal mulr_4_716 : std_logic_vector(9 downto 0);
    signal mulr_1_717 : std_logic_vector(9 downto 0);
    signal mulr_2_717 : std_logic_vector(9 downto 0);
    signal mulr_3_717 : std_logic_vector(9 downto 0);
    signal mulr_4_717 : std_logic_vector(9 downto 0);
    signal mulr_1_718 : std_logic_vector(9 downto 0);
    signal mulr_2_718 : std_logic_vector(9 downto 0);
    signal mulr_3_718 : std_logic_vector(9 downto 0);
    signal mulr_4_718 : std_logic_vector(9 downto 0);
    signal mulr_1_719 : std_logic_vector(9 downto 0);
    signal mulr_2_719 : std_logic_vector(9 downto 0);
    signal mulr_3_719 : std_logic_vector(9 downto 0);
    signal mulr_4_719 : std_logic_vector(9 downto 0);
    signal mulr_1_720 : std_logic_vector(9 downto 0);
    signal mulr_2_720 : std_logic_vector(9 downto 0);
    signal mulr_3_720 : std_logic_vector(9 downto 0);
    signal mulr_4_720 : std_logic_vector(9 downto 0);
    signal mulr_1_721 : std_logic_vector(9 downto 0);
    signal mulr_2_721 : std_logic_vector(9 downto 0);
    signal mulr_3_721 : std_logic_vector(9 downto 0);
    signal mulr_4_721 : std_logic_vector(9 downto 0);
    signal mulr_1_722 : std_logic_vector(9 downto 0);
    signal mulr_2_722 : std_logic_vector(9 downto 0);
    signal mulr_3_722 : std_logic_vector(9 downto 0);
    signal mulr_4_722 : std_logic_vector(9 downto 0);
    signal mulr_1_723 : std_logic_vector(9 downto 0);
    signal mulr_2_723 : std_logic_vector(9 downto 0);
    signal mulr_3_723 : std_logic_vector(9 downto 0);
    signal mulr_4_723 : std_logic_vector(9 downto 0);
    signal mulr_1_724 : std_logic_vector(9 downto 0);
    signal mulr_2_724 : std_logic_vector(9 downto 0);
    signal mulr_3_724 : std_logic_vector(9 downto 0);
    signal mulr_4_724 : std_logic_vector(9 downto 0);
    signal mulr_1_725 : std_logic_vector(9 downto 0);
    signal mulr_2_725 : std_logic_vector(9 downto 0);
    signal mulr_3_725 : std_logic_vector(9 downto 0);
    signal mulr_4_725 : std_logic_vector(9 downto 0);
    signal mulr_1_726 : std_logic_vector(9 downto 0);
    signal mulr_2_726 : std_logic_vector(9 downto 0);
    signal mulr_3_726 : std_logic_vector(9 downto 0);
    signal mulr_4_726 : std_logic_vector(9 downto 0);
    signal mulr_1_727 : std_logic_vector(9 downto 0);
    signal mulr_2_727 : std_logic_vector(9 downto 0);
    signal mulr_3_727 : std_logic_vector(9 downto 0);
    signal mulr_4_727 : std_logic_vector(9 downto 0);
    signal mulr_1_728 : std_logic_vector(9 downto 0);
    signal mulr_2_728 : std_logic_vector(9 downto 0);
    signal mulr_3_728 : std_logic_vector(9 downto 0);
    signal mulr_4_728 : std_logic_vector(9 downto 0);
    signal mulr_1_729 : std_logic_vector(9 downto 0);
    signal mulr_2_729 : std_logic_vector(9 downto 0);
    signal mulr_3_729 : std_logic_vector(9 downto 0);
    signal mulr_4_729 : std_logic_vector(9 downto 0);
    signal mulr_1_730 : std_logic_vector(9 downto 0);
    signal mulr_2_730 : std_logic_vector(9 downto 0);
    signal mulr_3_730 : std_logic_vector(9 downto 0);
    signal mulr_4_730 : std_logic_vector(9 downto 0);
    signal mulr_1_731 : std_logic_vector(9 downto 0);
    signal mulr_2_731 : std_logic_vector(9 downto 0);
    signal mulr_3_731 : std_logic_vector(9 downto 0);
    signal mulr_4_731 : std_logic_vector(9 downto 0);
    signal mulr_1_732 : std_logic_vector(9 downto 0);
    signal mulr_2_732 : std_logic_vector(9 downto 0);
    signal mulr_3_732 : std_logic_vector(9 downto 0);
    signal mulr_4_732 : std_logic_vector(9 downto 0);
    signal mulr_1_733 : std_logic_vector(9 downto 0);
    signal mulr_2_733 : std_logic_vector(9 downto 0);
    signal mulr_3_733 : std_logic_vector(9 downto 0);
    signal mulr_4_733 : std_logic_vector(9 downto 0);
    signal mulr_1_734 : std_logic_vector(9 downto 0);
    signal mulr_2_734 : std_logic_vector(9 downto 0);
    signal mulr_3_734 : std_logic_vector(9 downto 0);
    signal mulr_4_734 : std_logic_vector(9 downto 0);
    signal mulr_1_735 : std_logic_vector(9 downto 0);
    signal mulr_2_735 : std_logic_vector(9 downto 0);
    signal mulr_3_735 : std_logic_vector(9 downto 0);
    signal mulr_4_735 : std_logic_vector(9 downto 0);
    signal mulr_1_736 : std_logic_vector(9 downto 0);
    signal mulr_2_736 : std_logic_vector(9 downto 0);
    signal mulr_3_736 : std_logic_vector(9 downto 0);
    signal mulr_4_736 : std_logic_vector(9 downto 0);
    signal mulr_1_737 : std_logic_vector(9 downto 0);
    signal mulr_2_737 : std_logic_vector(9 downto 0);
    signal mulr_3_737 : std_logic_vector(9 downto 0);
    signal mulr_4_737 : std_logic_vector(9 downto 0);
    signal mulr_1_738 : std_logic_vector(9 downto 0);
    signal mulr_2_738 : std_logic_vector(9 downto 0);
    signal mulr_3_738 : std_logic_vector(9 downto 0);
    signal mulr_4_738 : std_logic_vector(9 downto 0);
    signal mulr_1_739 : std_logic_vector(9 downto 0);
    signal mulr_2_739 : std_logic_vector(9 downto 0);
    signal mulr_3_739 : std_logic_vector(9 downto 0);
    signal mulr_4_739 : std_logic_vector(9 downto 0);
    signal mulr_1_740 : std_logic_vector(9 downto 0);
    signal mulr_2_740 : std_logic_vector(9 downto 0);
    signal mulr_3_740 : std_logic_vector(9 downto 0);
    signal mulr_4_740 : std_logic_vector(9 downto 0);
    signal mulr_1_741 : std_logic_vector(9 downto 0);
    signal mulr_2_741 : std_logic_vector(9 downto 0);
    signal mulr_3_741 : std_logic_vector(9 downto 0);
    signal mulr_4_741 : std_logic_vector(9 downto 0);
    signal mulr_1_742 : std_logic_vector(9 downto 0);
    signal mulr_2_742 : std_logic_vector(9 downto 0);
    signal mulr_3_742 : std_logic_vector(9 downto 0);
    signal mulr_4_742 : std_logic_vector(9 downto 0);
    signal mulr_1_743 : std_logic_vector(9 downto 0);
    signal mulr_2_743 : std_logic_vector(9 downto 0);
    signal mulr_3_743 : std_logic_vector(9 downto 0);
    signal mulr_4_743 : std_logic_vector(9 downto 0);
    signal mulr_1_744 : std_logic_vector(9 downto 0);
    signal mulr_2_744 : std_logic_vector(9 downto 0);
    signal mulr_3_744 : std_logic_vector(9 downto 0);
    signal mulr_4_744 : std_logic_vector(9 downto 0);
    signal mulr_1_745 : std_logic_vector(9 downto 0);
    signal mulr_2_745 : std_logic_vector(9 downto 0);
    signal mulr_3_745 : std_logic_vector(9 downto 0);
    signal mulr_4_745 : std_logic_vector(9 downto 0);
    signal mulr_1_746 : std_logic_vector(9 downto 0);
    signal mulr_2_746 : std_logic_vector(9 downto 0);
    signal mulr_3_746 : std_logic_vector(9 downto 0);
    signal mulr_4_746 : std_logic_vector(9 downto 0);
    signal mulr_1_747 : std_logic_vector(9 downto 0);
    signal mulr_2_747 : std_logic_vector(9 downto 0);
    signal mulr_3_747 : std_logic_vector(9 downto 0);
    signal mulr_4_747 : std_logic_vector(9 downto 0);
    signal mulr_1_748 : std_logic_vector(9 downto 0);
    signal mulr_2_748 : std_logic_vector(9 downto 0);
    signal mulr_3_748 : std_logic_vector(9 downto 0);
    signal mulr_4_748 : std_logic_vector(9 downto 0);
    signal mulr_1_749 : std_logic_vector(9 downto 0);
    signal mulr_2_749 : std_logic_vector(9 downto 0);
    signal mulr_3_749 : std_logic_vector(9 downto 0);
    signal mulr_4_749 : std_logic_vector(9 downto 0);
    signal mulr_1_750 : std_logic_vector(9 downto 0);
    signal mulr_2_750 : std_logic_vector(9 downto 0);
    signal mulr_3_750 : std_logic_vector(9 downto 0);
    signal mulr_4_750 : std_logic_vector(9 downto 0);
    signal mulr_1_751 : std_logic_vector(9 downto 0);
    signal mulr_2_751 : std_logic_vector(9 downto 0);
    signal mulr_3_751 : std_logic_vector(9 downto 0);
    signal mulr_4_751 : std_logic_vector(9 downto 0);
    signal mulr_1_752 : std_logic_vector(9 downto 0);
    signal mulr_2_752 : std_logic_vector(9 downto 0);
    signal mulr_3_752 : std_logic_vector(9 downto 0);
    signal mulr_4_752 : std_logic_vector(9 downto 0);
    signal mulr_1_753 : std_logic_vector(9 downto 0);
    signal mulr_2_753 : std_logic_vector(9 downto 0);
    signal mulr_3_753 : std_logic_vector(9 downto 0);
    signal mulr_4_753 : std_logic_vector(9 downto 0);
    signal mulr_1_754 : std_logic_vector(9 downto 0);
    signal mulr_2_754 : std_logic_vector(9 downto 0);
    signal mulr_3_754 : std_logic_vector(9 downto 0);
    signal mulr_4_754 : std_logic_vector(9 downto 0);
    signal mulr_1_755 : std_logic_vector(9 downto 0);
    signal mulr_2_755 : std_logic_vector(9 downto 0);
    signal mulr_3_755 : std_logic_vector(9 downto 0);
    signal mulr_4_755 : std_logic_vector(9 downto 0);
    signal mulr_1_756 : std_logic_vector(9 downto 0);
    signal mulr_2_756 : std_logic_vector(9 downto 0);
    signal mulr_3_756 : std_logic_vector(9 downto 0);
    signal mulr_4_756 : std_logic_vector(9 downto 0);
    signal mulr_1_757 : std_logic_vector(9 downto 0);
    signal mulr_2_757 : std_logic_vector(9 downto 0);
    signal mulr_3_757 : std_logic_vector(9 downto 0);
    signal mulr_4_757 : std_logic_vector(9 downto 0);
    signal mulr_1_758 : std_logic_vector(9 downto 0);
    signal mulr_2_758 : std_logic_vector(9 downto 0);
    signal mulr_3_758 : std_logic_vector(9 downto 0);
    signal mulr_4_758 : std_logic_vector(9 downto 0);
    signal mulr_1_759 : std_logic_vector(9 downto 0);
    signal mulr_2_759 : std_logic_vector(9 downto 0);
    signal mulr_3_759 : std_logic_vector(9 downto 0);
    signal mulr_4_759 : std_logic_vector(9 downto 0);
    signal mulr_1_760 : std_logic_vector(9 downto 0);
    signal mulr_2_760 : std_logic_vector(9 downto 0);
    signal mulr_3_760 : std_logic_vector(9 downto 0);
    signal mulr_4_760 : std_logic_vector(9 downto 0);
    signal mulr_1_761 : std_logic_vector(9 downto 0);
    signal mulr_2_761 : std_logic_vector(9 downto 0);
    signal mulr_3_761 : std_logic_vector(9 downto 0);
    signal mulr_4_761 : std_logic_vector(9 downto 0);
    signal mulr_1_762 : std_logic_vector(9 downto 0);
    signal mulr_2_762 : std_logic_vector(9 downto 0);
    signal mulr_3_762 : std_logic_vector(9 downto 0);
    signal mulr_4_762 : std_logic_vector(9 downto 0);
    signal mulr_1_763 : std_logic_vector(9 downto 0);
    signal mulr_2_763 : std_logic_vector(9 downto 0);
    signal mulr_3_763 : std_logic_vector(9 downto 0);
    signal mulr_4_763 : std_logic_vector(9 downto 0);
    signal mulr_1_764 : std_logic_vector(9 downto 0);
    signal mulr_2_764 : std_logic_vector(9 downto 0);
    signal mulr_3_764 : std_logic_vector(9 downto 0);
    signal mulr_4_764 : std_logic_vector(9 downto 0);
    signal mulr_1_765 : std_logic_vector(9 downto 0);
    signal mulr_2_765 : std_logic_vector(9 downto 0);
    signal mulr_3_765 : std_logic_vector(9 downto 0);
    signal mulr_4_765 : std_logic_vector(9 downto 0);
    signal mulr_1_766 : std_logic_vector(9 downto 0);
    signal mulr_2_766 : std_logic_vector(9 downto 0);
    signal mulr_3_766 : std_logic_vector(9 downto 0);
    signal mulr_4_766 : std_logic_vector(9 downto 0);
    signal mulr_1_767 : std_logic_vector(9 downto 0);
    signal mulr_2_767 : std_logic_vector(9 downto 0);
    signal mulr_3_767 : std_logic_vector(9 downto 0);
    signal mulr_4_767 : std_logic_vector(9 downto 0);
    signal mulr_1_768 : std_logic_vector(9 downto 0);
    signal mulr_2_768 : std_logic_vector(9 downto 0);
    signal mulr_3_768 : std_logic_vector(9 downto 0);
    signal mulr_4_768 : std_logic_vector(9 downto 0);
    signal mulr_1_769 : std_logic_vector(9 downto 0);
    signal mulr_2_769 : std_logic_vector(9 downto 0);
    signal mulr_3_769 : std_logic_vector(9 downto 0);
    signal mulr_4_769 : std_logic_vector(9 downto 0);
    signal mulr_1_770 : std_logic_vector(9 downto 0);
    signal mulr_2_770 : std_logic_vector(9 downto 0);
    signal mulr_3_770 : std_logic_vector(9 downto 0);
    signal mulr_4_770 : std_logic_vector(9 downto 0);
    signal mulr_1_771 : std_logic_vector(9 downto 0);
    signal mulr_2_771 : std_logic_vector(9 downto 0);
    signal mulr_3_771 : std_logic_vector(9 downto 0);
    signal mulr_4_771 : std_logic_vector(9 downto 0);
    signal mulr_1_772 : std_logic_vector(9 downto 0);
    signal mulr_2_772 : std_logic_vector(9 downto 0);
    signal mulr_3_772 : std_logic_vector(9 downto 0);
    signal mulr_4_772 : std_logic_vector(9 downto 0);
    signal mulr_1_773 : std_logic_vector(9 downto 0);
    signal mulr_2_773 : std_logic_vector(9 downto 0);
    signal mulr_3_773 : std_logic_vector(9 downto 0);
    signal mulr_4_773 : std_logic_vector(9 downto 0);
    signal mulr_1_774 : std_logic_vector(9 downto 0);
    signal mulr_2_774 : std_logic_vector(9 downto 0);
    signal mulr_3_774 : std_logic_vector(9 downto 0);
    signal mulr_4_774 : std_logic_vector(9 downto 0);
    signal mulr_1_775 : std_logic_vector(9 downto 0);
    signal mulr_2_775 : std_logic_vector(9 downto 0);
    signal mulr_3_775 : std_logic_vector(9 downto 0);
    signal mulr_4_775 : std_logic_vector(9 downto 0);
    signal mulr_1_776 : std_logic_vector(9 downto 0);
    signal mulr_2_776 : std_logic_vector(9 downto 0);
    signal mulr_3_776 : std_logic_vector(9 downto 0);
    signal mulr_4_776 : std_logic_vector(9 downto 0);
    signal mulr_1_777 : std_logic_vector(9 downto 0);
    signal mulr_2_777 : std_logic_vector(9 downto 0);
    signal mulr_3_777 : std_logic_vector(9 downto 0);
    signal mulr_4_777 : std_logic_vector(9 downto 0);
    signal mulr_1_778 : std_logic_vector(9 downto 0);
    signal mulr_2_778 : std_logic_vector(9 downto 0);
    signal mulr_3_778 : std_logic_vector(9 downto 0);
    signal mulr_4_778 : std_logic_vector(9 downto 0);
    signal mulr_1_779 : std_logic_vector(9 downto 0);
    signal mulr_2_779 : std_logic_vector(9 downto 0);
    signal mulr_3_779 : std_logic_vector(9 downto 0);
    signal mulr_4_779 : std_logic_vector(9 downto 0);
    signal mulr_1_780 : std_logic_vector(9 downto 0);
    signal mulr_2_780 : std_logic_vector(9 downto 0);
    signal mulr_3_780 : std_logic_vector(9 downto 0);
    signal mulr_4_780 : std_logic_vector(9 downto 0);
    signal mulr_1_781 : std_logic_vector(9 downto 0);
    signal mulr_2_781 : std_logic_vector(9 downto 0);
    signal mulr_3_781 : std_logic_vector(9 downto 0);
    signal mulr_4_781 : std_logic_vector(9 downto 0);
    signal mulr_1_782 : std_logic_vector(9 downto 0);
    signal mulr_2_782 : std_logic_vector(9 downto 0);
    signal mulr_3_782 : std_logic_vector(9 downto 0);
    signal mulr_4_782 : std_logic_vector(9 downto 0);
    signal mulr_1_783 : std_logic_vector(9 downto 0);
    signal mulr_2_783 : std_logic_vector(9 downto 0);
    signal mulr_3_783 : std_logic_vector(9 downto 0);
    signal mulr_4_783 : std_logic_vector(9 downto 0);
    signal mulr_1_784 : std_logic_vector(9 downto 0);
    signal mulr_2_784 : std_logic_vector(9 downto 0);
    signal mulr_3_784 : std_logic_vector(9 downto 0);
    signal mulr_4_784 : std_logic_vector(9 downto 0);
    signal mulr_1_785 : std_logic_vector(9 downto 0);
    signal mulr_2_785 : std_logic_vector(9 downto 0);
    signal mulr_3_785 : std_logic_vector(9 downto 0);
    signal mulr_4_785 : std_logic_vector(9 downto 0);
    signal mulr_1_786 : std_logic_vector(9 downto 0);
    signal mulr_2_786 : std_logic_vector(9 downto 0);
    signal mulr_3_786 : std_logic_vector(9 downto 0);
    signal mulr_4_786 : std_logic_vector(9 downto 0);
    signal mulr_1_787 : std_logic_vector(9 downto 0);
    signal mulr_2_787 : std_logic_vector(9 downto 0);
    signal mulr_3_787 : std_logic_vector(9 downto 0);
    signal mulr_4_787 : std_logic_vector(9 downto 0);
    signal mulr_1_788 : std_logic_vector(9 downto 0);
    signal mulr_2_788 : std_logic_vector(9 downto 0);
    signal mulr_3_788 : std_logic_vector(9 downto 0);
    signal mulr_4_788 : std_logic_vector(9 downto 0);
    signal mulr_1_789 : std_logic_vector(9 downto 0);
    signal mulr_2_789 : std_logic_vector(9 downto 0);
    signal mulr_3_789 : std_logic_vector(9 downto 0);
    signal mulr_4_789 : std_logic_vector(9 downto 0);
    signal mulr_1_790 : std_logic_vector(9 downto 0);
    signal mulr_2_790 : std_logic_vector(9 downto 0);
    signal mulr_3_790 : std_logic_vector(9 downto 0);
    signal mulr_4_790 : std_logic_vector(9 downto 0);
    signal mulr_1_791 : std_logic_vector(9 downto 0);
    signal mulr_2_791 : std_logic_vector(9 downto 0);
    signal mulr_3_791 : std_logic_vector(9 downto 0);
    signal mulr_4_791 : std_logic_vector(9 downto 0);
    signal mulr_1_792 : std_logic_vector(9 downto 0);
    signal mulr_2_792 : std_logic_vector(9 downto 0);
    signal mulr_3_792 : std_logic_vector(9 downto 0);
    signal mulr_4_792 : std_logic_vector(9 downto 0);
    signal mulr_1_793 : std_logic_vector(9 downto 0);
    signal mulr_2_793 : std_logic_vector(9 downto 0);
    signal mulr_3_793 : std_logic_vector(9 downto 0);
    signal mulr_4_793 : std_logic_vector(9 downto 0);
    signal mulr_1_794 : std_logic_vector(9 downto 0);
    signal mulr_2_794 : std_logic_vector(9 downto 0);
    signal mulr_3_794 : std_logic_vector(9 downto 0);
    signal mulr_4_794 : std_logic_vector(9 downto 0);
    signal mulr_1_795 : std_logic_vector(9 downto 0);
    signal mulr_2_795 : std_logic_vector(9 downto 0);
    signal mulr_3_795 : std_logic_vector(9 downto 0);
    signal mulr_4_795 : std_logic_vector(9 downto 0);
    signal mulr_1_796 : std_logic_vector(9 downto 0);
    signal mulr_2_796 : std_logic_vector(9 downto 0);
    signal mulr_3_796 : std_logic_vector(9 downto 0);
    signal mulr_4_796 : std_logic_vector(9 downto 0);
    signal mulr_1_797 : std_logic_vector(9 downto 0);
    signal mulr_2_797 : std_logic_vector(9 downto 0);
    signal mulr_3_797 : std_logic_vector(9 downto 0);
    signal mulr_4_797 : std_logic_vector(9 downto 0);
    signal mulr_1_798 : std_logic_vector(9 downto 0);
    signal mulr_2_798 : std_logic_vector(9 downto 0);
    signal mulr_3_798 : std_logic_vector(9 downto 0);
    signal mulr_4_798 : std_logic_vector(9 downto 0);
    signal mulr_1_799 : std_logic_vector(9 downto 0);
    signal mulr_2_799 : std_logic_vector(9 downto 0);
    signal mulr_3_799 : std_logic_vector(9 downto 0);
    signal mulr_4_799 : std_logic_vector(9 downto 0);
    signal mulr_1_800 : std_logic_vector(9 downto 0);
    signal mulr_2_800 : std_logic_vector(9 downto 0);
    signal mulr_3_800 : std_logic_vector(9 downto 0);
    signal mulr_4_800 : std_logic_vector(9 downto 0);
    signal mulr_1_801 : std_logic_vector(9 downto 0);
    signal mulr_2_801 : std_logic_vector(9 downto 0);
    signal mulr_3_801 : std_logic_vector(9 downto 0);
    signal mulr_4_801 : std_logic_vector(9 downto 0);
    signal mulr_1_802 : std_logic_vector(9 downto 0);
    signal mulr_2_802 : std_logic_vector(9 downto 0);
    signal mulr_3_802 : std_logic_vector(9 downto 0);
    signal mulr_4_802 : std_logic_vector(9 downto 0);
    signal mulr_1_803 : std_logic_vector(9 downto 0);
    signal mulr_2_803 : std_logic_vector(9 downto 0);
    signal mulr_3_803 : std_logic_vector(9 downto 0);
    signal mulr_4_803 : std_logic_vector(9 downto 0);
    signal mulr_1_804 : std_logic_vector(9 downto 0);
    signal mulr_2_804 : std_logic_vector(9 downto 0);
    signal mulr_3_804 : std_logic_vector(9 downto 0);
    signal mulr_4_804 : std_logic_vector(9 downto 0);
    signal mulr_1_805 : std_logic_vector(9 downto 0);
    signal mulr_2_805 : std_logic_vector(9 downto 0);
    signal mulr_3_805 : std_logic_vector(9 downto 0);
    signal mulr_4_805 : std_logic_vector(9 downto 0);
    signal mulr_1_806 : std_logic_vector(9 downto 0);
    signal mulr_2_806 : std_logic_vector(9 downto 0);
    signal mulr_3_806 : std_logic_vector(9 downto 0);
    signal mulr_4_806 : std_logic_vector(9 downto 0);
    signal mulr_1_807 : std_logic_vector(9 downto 0);
    signal mulr_2_807 : std_logic_vector(9 downto 0);
    signal mulr_3_807 : std_logic_vector(9 downto 0);
    signal mulr_4_807 : std_logic_vector(9 downto 0);
    signal mulr_1_808 : std_logic_vector(9 downto 0);
    signal mulr_2_808 : std_logic_vector(9 downto 0);
    signal mulr_3_808 : std_logic_vector(9 downto 0);
    signal mulr_4_808 : std_logic_vector(9 downto 0);
    signal mulr_1_809 : std_logic_vector(9 downto 0);
    signal mulr_2_809 : std_logic_vector(9 downto 0);
    signal mulr_3_809 : std_logic_vector(9 downto 0);
    signal mulr_4_809 : std_logic_vector(9 downto 0);
    signal mulr_1_810 : std_logic_vector(9 downto 0);
    signal mulr_2_810 : std_logic_vector(9 downto 0);
    signal mulr_3_810 : std_logic_vector(9 downto 0);
    signal mulr_4_810 : std_logic_vector(9 downto 0);
    signal mulr_1_811 : std_logic_vector(9 downto 0);
    signal mulr_2_811 : std_logic_vector(9 downto 0);
    signal mulr_3_811 : std_logic_vector(9 downto 0);
    signal mulr_4_811 : std_logic_vector(9 downto 0);
    signal mulr_1_812 : std_logic_vector(9 downto 0);
    signal mulr_2_812 : std_logic_vector(9 downto 0);
    signal mulr_3_812 : std_logic_vector(9 downto 0);
    signal mulr_4_812 : std_logic_vector(9 downto 0);
    signal mulr_1_813 : std_logic_vector(9 downto 0);
    signal mulr_2_813 : std_logic_vector(9 downto 0);
    signal mulr_3_813 : std_logic_vector(9 downto 0);
    signal mulr_4_813 : std_logic_vector(9 downto 0);
    signal mulr_1_814 : std_logic_vector(9 downto 0);
    signal mulr_2_814 : std_logic_vector(9 downto 0);
    signal mulr_3_814 : std_logic_vector(9 downto 0);
    signal mulr_4_814 : std_logic_vector(9 downto 0);
    signal mulr_1_815 : std_logic_vector(9 downto 0);
    signal mulr_2_815 : std_logic_vector(9 downto 0);
    signal mulr_3_815 : std_logic_vector(9 downto 0);
    signal mulr_4_815 : std_logic_vector(9 downto 0);
    signal mulr_1_816 : std_logic_vector(9 downto 0);
    signal mulr_2_816 : std_logic_vector(9 downto 0);
    signal mulr_3_816 : std_logic_vector(9 downto 0);
    signal mulr_4_816 : std_logic_vector(9 downto 0);
    signal mulr_1_817 : std_logic_vector(9 downto 0);
    signal mulr_2_817 : std_logic_vector(9 downto 0);
    signal mulr_3_817 : std_logic_vector(9 downto 0);
    signal mulr_4_817 : std_logic_vector(9 downto 0);
    signal mulr_1_818 : std_logic_vector(9 downto 0);
    signal mulr_2_818 : std_logic_vector(9 downto 0);
    signal mulr_3_818 : std_logic_vector(9 downto 0);
    signal mulr_4_818 : std_logic_vector(9 downto 0);
    signal mulr_1_819 : std_logic_vector(9 downto 0);
    signal mulr_2_819 : std_logic_vector(9 downto 0);
    signal mulr_3_819 : std_logic_vector(9 downto 0);
    signal mulr_4_819 : std_logic_vector(9 downto 0);
    signal mulr_1_820 : std_logic_vector(9 downto 0);
    signal mulr_2_820 : std_logic_vector(9 downto 0);
    signal mulr_3_820 : std_logic_vector(9 downto 0);
    signal mulr_4_820 : std_logic_vector(9 downto 0);
    signal mulr_1_821 : std_logic_vector(9 downto 0);
    signal mulr_2_821 : std_logic_vector(9 downto 0);
    signal mulr_3_821 : std_logic_vector(9 downto 0);
    signal mulr_4_821 : std_logic_vector(9 downto 0);
    signal mulr_1_822 : std_logic_vector(9 downto 0);
    signal mulr_2_822 : std_logic_vector(9 downto 0);
    signal mulr_3_822 : std_logic_vector(9 downto 0);
    signal mulr_4_822 : std_logic_vector(9 downto 0);
    signal mulr_1_823 : std_logic_vector(9 downto 0);
    signal mulr_2_823 : std_logic_vector(9 downto 0);
    signal mulr_3_823 : std_logic_vector(9 downto 0);
    signal mulr_4_823 : std_logic_vector(9 downto 0);
    signal mulr_1_824 : std_logic_vector(9 downto 0);
    signal mulr_2_824 : std_logic_vector(9 downto 0);
    signal mulr_3_824 : std_logic_vector(9 downto 0);
    signal mulr_4_824 : std_logic_vector(9 downto 0);
    signal mulr_1_825 : std_logic_vector(9 downto 0);
    signal mulr_2_825 : std_logic_vector(9 downto 0);
    signal mulr_3_825 : std_logic_vector(9 downto 0);
    signal mulr_4_825 : std_logic_vector(9 downto 0);
    signal mulr_1_826 : std_logic_vector(9 downto 0);
    signal mulr_2_826 : std_logic_vector(9 downto 0);
    signal mulr_3_826 : std_logic_vector(9 downto 0);
    signal mulr_4_826 : std_logic_vector(9 downto 0);
    signal mulr_1_827 : std_logic_vector(9 downto 0);
    signal mulr_2_827 : std_logic_vector(9 downto 0);
    signal mulr_3_827 : std_logic_vector(9 downto 0);
    signal mulr_4_827 : std_logic_vector(9 downto 0);
    signal mulr_1_828 : std_logic_vector(9 downto 0);
    signal mulr_2_828 : std_logic_vector(9 downto 0);
    signal mulr_3_828 : std_logic_vector(9 downto 0);
    signal mulr_4_828 : std_logic_vector(9 downto 0);
    signal mulr_1_829 : std_logic_vector(9 downto 0);
    signal mulr_2_829 : std_logic_vector(9 downto 0);
    signal mulr_3_829 : std_logic_vector(9 downto 0);
    signal mulr_4_829 : std_logic_vector(9 downto 0);
    signal mulr_1_830 : std_logic_vector(9 downto 0);
    signal mulr_2_830 : std_logic_vector(9 downto 0);
    signal mulr_3_830 : std_logic_vector(9 downto 0);
    signal mulr_4_830 : std_logic_vector(9 downto 0);
    signal mulr_1_831 : std_logic_vector(9 downto 0);
    signal mulr_2_831 : std_logic_vector(9 downto 0);
    signal mulr_3_831 : std_logic_vector(9 downto 0);
    signal mulr_4_831 : std_logic_vector(9 downto 0);
    signal mulr_1_832 : std_logic_vector(9 downto 0);
    signal mulr_2_832 : std_logic_vector(9 downto 0);
    signal mulr_3_832 : std_logic_vector(9 downto 0);
    signal mulr_4_832 : std_logic_vector(9 downto 0);
    signal mulr_1_833 : std_logic_vector(9 downto 0);
    signal mulr_2_833 : std_logic_vector(9 downto 0);
    signal mulr_3_833 : std_logic_vector(9 downto 0);
    signal mulr_4_833 : std_logic_vector(9 downto 0);
    signal mulr_1_834 : std_logic_vector(9 downto 0);
    signal mulr_2_834 : std_logic_vector(9 downto 0);
    signal mulr_3_834 : std_logic_vector(9 downto 0);
    signal mulr_4_834 : std_logic_vector(9 downto 0);
    signal mulr_1_835 : std_logic_vector(9 downto 0);
    signal mulr_2_835 : std_logic_vector(9 downto 0);
    signal mulr_3_835 : std_logic_vector(9 downto 0);
    signal mulr_4_835 : std_logic_vector(9 downto 0);
    signal mulr_1_836 : std_logic_vector(9 downto 0);
    signal mulr_2_836 : std_logic_vector(9 downto 0);
    signal mulr_3_836 : std_logic_vector(9 downto 0);
    signal mulr_4_836 : std_logic_vector(9 downto 0);
    signal mulr_1_837 : std_logic_vector(9 downto 0);
    signal mulr_2_837 : std_logic_vector(9 downto 0);
    signal mulr_3_837 : std_logic_vector(9 downto 0);
    signal mulr_4_837 : std_logic_vector(9 downto 0);
    signal mulr_1_838 : std_logic_vector(9 downto 0);
    signal mulr_2_838 : std_logic_vector(9 downto 0);
    signal mulr_3_838 : std_logic_vector(9 downto 0);
    signal mulr_4_838 : std_logic_vector(9 downto 0);
    signal mulr_1_839 : std_logic_vector(9 downto 0);
    signal mulr_2_839 : std_logic_vector(9 downto 0);
    signal mulr_3_839 : std_logic_vector(9 downto 0);
    signal mulr_4_839 : std_logic_vector(9 downto 0);
    signal mulr_1_840 : std_logic_vector(9 downto 0);
    signal mulr_2_840 : std_logic_vector(9 downto 0);
    signal mulr_3_840 : std_logic_vector(9 downto 0);
    signal mulr_4_840 : std_logic_vector(9 downto 0);
    signal mulr_1_841 : std_logic_vector(9 downto 0);
    signal mulr_2_841 : std_logic_vector(9 downto 0);
    signal mulr_3_841 : std_logic_vector(9 downto 0);
    signal mulr_4_841 : std_logic_vector(9 downto 0);
    signal mulr_1_842 : std_logic_vector(9 downto 0);
    signal mulr_2_842 : std_logic_vector(9 downto 0);
    signal mulr_3_842 : std_logic_vector(9 downto 0);
    signal mulr_4_842 : std_logic_vector(9 downto 0);
    signal mulr_1_843 : std_logic_vector(9 downto 0);
    signal mulr_2_843 : std_logic_vector(9 downto 0);
    signal mulr_3_843 : std_logic_vector(9 downto 0);
    signal mulr_4_843 : std_logic_vector(9 downto 0);
    signal mulr_1_844 : std_logic_vector(9 downto 0);
    signal mulr_2_844 : std_logic_vector(9 downto 0);
    signal mulr_3_844 : std_logic_vector(9 downto 0);
    signal mulr_4_844 : std_logic_vector(9 downto 0);
    signal mulr_1_845 : std_logic_vector(9 downto 0);
    signal mulr_2_845 : std_logic_vector(9 downto 0);
    signal mulr_3_845 : std_logic_vector(9 downto 0);
    signal mulr_4_845 : std_logic_vector(9 downto 0);
    signal mulr_1_846 : std_logic_vector(9 downto 0);
    signal mulr_2_846 : std_logic_vector(9 downto 0);
    signal mulr_3_846 : std_logic_vector(9 downto 0);
    signal mulr_4_846 : std_logic_vector(9 downto 0);
    signal mulr_1_847 : std_logic_vector(9 downto 0);
    signal mulr_2_847 : std_logic_vector(9 downto 0);
    signal mulr_3_847 : std_logic_vector(9 downto 0);
    signal mulr_4_847 : std_logic_vector(9 downto 0);
    signal mulr_1_848 : std_logic_vector(9 downto 0);
    signal mulr_2_848 : std_logic_vector(9 downto 0);
    signal mulr_3_848 : std_logic_vector(9 downto 0);
    signal mulr_4_848 : std_logic_vector(9 downto 0);
    signal mulr_1_849 : std_logic_vector(9 downto 0);
    signal mulr_2_849 : std_logic_vector(9 downto 0);
    signal mulr_3_849 : std_logic_vector(9 downto 0);
    signal mulr_4_849 : std_logic_vector(9 downto 0);
    signal mulr_1_850 : std_logic_vector(9 downto 0);
    signal mulr_2_850 : std_logic_vector(9 downto 0);
    signal mulr_3_850 : std_logic_vector(9 downto 0);
    signal mulr_4_850 : std_logic_vector(9 downto 0);
    signal mulr_1_851 : std_logic_vector(9 downto 0);
    signal mulr_2_851 : std_logic_vector(9 downto 0);
    signal mulr_3_851 : std_logic_vector(9 downto 0);
    signal mulr_4_851 : std_logic_vector(9 downto 0);
    signal mulr_1_852 : std_logic_vector(9 downto 0);
    signal mulr_2_852 : std_logic_vector(9 downto 0);
    signal mulr_3_852 : std_logic_vector(9 downto 0);
    signal mulr_4_852 : std_logic_vector(9 downto 0);
    signal mulr_1_853 : std_logic_vector(9 downto 0);
    signal mulr_2_853 : std_logic_vector(9 downto 0);
    signal mulr_3_853 : std_logic_vector(9 downto 0);
    signal mulr_4_853 : std_logic_vector(9 downto 0);
    signal mulr_1_854 : std_logic_vector(9 downto 0);
    signal mulr_2_854 : std_logic_vector(9 downto 0);
    signal mulr_3_854 : std_logic_vector(9 downto 0);
    signal mulr_4_854 : std_logic_vector(9 downto 0);
    signal mulr_1_855 : std_logic_vector(9 downto 0);
    signal mulr_2_855 : std_logic_vector(9 downto 0);
    signal mulr_3_855 : std_logic_vector(9 downto 0);
    signal mulr_4_855 : std_logic_vector(9 downto 0);
    signal mulr_1_856 : std_logic_vector(9 downto 0);
    signal mulr_2_856 : std_logic_vector(9 downto 0);
    signal mulr_3_856 : std_logic_vector(9 downto 0);
    signal mulr_4_856 : std_logic_vector(9 downto 0);
    signal mulr_1_857 : std_logic_vector(9 downto 0);
    signal mulr_2_857 : std_logic_vector(9 downto 0);
    signal mulr_3_857 : std_logic_vector(9 downto 0);
    signal mulr_4_857 : std_logic_vector(9 downto 0);
    signal mulr_1_858 : std_logic_vector(9 downto 0);
    signal mulr_2_858 : std_logic_vector(9 downto 0);
    signal mulr_3_858 : std_logic_vector(9 downto 0);
    signal mulr_4_858 : std_logic_vector(9 downto 0);
    signal mulr_1_859 : std_logic_vector(9 downto 0);
    signal mulr_2_859 : std_logic_vector(9 downto 0);
    signal mulr_3_859 : std_logic_vector(9 downto 0);
    signal mulr_4_859 : std_logic_vector(9 downto 0);
    signal mulr_1_860 : std_logic_vector(9 downto 0);
    signal mulr_2_860 : std_logic_vector(9 downto 0);
    signal mulr_3_860 : std_logic_vector(9 downto 0);
    signal mulr_4_860 : std_logic_vector(9 downto 0);
    signal mulr_1_861 : std_logic_vector(9 downto 0);
    signal mulr_2_861 : std_logic_vector(9 downto 0);
    signal mulr_3_861 : std_logic_vector(9 downto 0);
    signal mulr_4_861 : std_logic_vector(9 downto 0);
    signal mulr_1_862 : std_logic_vector(9 downto 0);
    signal mulr_2_862 : std_logic_vector(9 downto 0);
    signal mulr_3_862 : std_logic_vector(9 downto 0);
    signal mulr_4_862 : std_logic_vector(9 downto 0);
    signal mulr_1_863 : std_logic_vector(9 downto 0);
    signal mulr_2_863 : std_logic_vector(9 downto 0);
    signal mulr_3_863 : std_logic_vector(9 downto 0);
    signal mulr_4_863 : std_logic_vector(9 downto 0);
    signal mulr_1_864 : std_logic_vector(9 downto 0);
    signal mulr_2_864 : std_logic_vector(9 downto 0);
    signal mulr_3_864 : std_logic_vector(9 downto 0);
    signal mulr_4_864 : std_logic_vector(9 downto 0);
    signal mulr_1_865 : std_logic_vector(9 downto 0);
    signal mulr_2_865 : std_logic_vector(9 downto 0);
    signal mulr_3_865 : std_logic_vector(9 downto 0);
    signal mulr_4_865 : std_logic_vector(9 downto 0);
    signal mulr_1_866 : std_logic_vector(9 downto 0);
    signal mulr_2_866 : std_logic_vector(9 downto 0);
    signal mulr_3_866 : std_logic_vector(9 downto 0);
    signal mulr_4_866 : std_logic_vector(9 downto 0);
    signal mulr_1_867 : std_logic_vector(9 downto 0);
    signal mulr_2_867 : std_logic_vector(9 downto 0);
    signal mulr_3_867 : std_logic_vector(9 downto 0);
    signal mulr_4_867 : std_logic_vector(9 downto 0);
    signal mulr_1_868 : std_logic_vector(9 downto 0);
    signal mulr_2_868 : std_logic_vector(9 downto 0);
    signal mulr_3_868 : std_logic_vector(9 downto 0);
    signal mulr_4_868 : std_logic_vector(9 downto 0);
    signal mulr_1_869 : std_logic_vector(9 downto 0);
    signal mulr_2_869 : std_logic_vector(9 downto 0);
    signal mulr_3_869 : std_logic_vector(9 downto 0);
    signal mulr_4_869 : std_logic_vector(9 downto 0);
    signal mulr_1_870 : std_logic_vector(9 downto 0);
    signal mulr_2_870 : std_logic_vector(9 downto 0);
    signal mulr_3_870 : std_logic_vector(9 downto 0);
    signal mulr_4_870 : std_logic_vector(9 downto 0);
    signal mulr_1_871 : std_logic_vector(9 downto 0);
    signal mulr_2_871 : std_logic_vector(9 downto 0);
    signal mulr_3_871 : std_logic_vector(9 downto 0);
    signal mulr_4_871 : std_logic_vector(9 downto 0);
    signal mulr_1_872 : std_logic_vector(9 downto 0);
    signal mulr_2_872 : std_logic_vector(9 downto 0);
    signal mulr_3_872 : std_logic_vector(9 downto 0);
    signal mulr_4_872 : std_logic_vector(9 downto 0);
    signal mulr_1_873 : std_logic_vector(9 downto 0);
    signal mulr_2_873 : std_logic_vector(9 downto 0);
    signal mulr_3_873 : std_logic_vector(9 downto 0);
    signal mulr_4_873 : std_logic_vector(9 downto 0);
    signal mulr_1_874 : std_logic_vector(9 downto 0);
    signal mulr_2_874 : std_logic_vector(9 downto 0);
    signal mulr_3_874 : std_logic_vector(9 downto 0);
    signal mulr_4_874 : std_logic_vector(9 downto 0);
    signal mulr_1_875 : std_logic_vector(9 downto 0);
    signal mulr_2_875 : std_logic_vector(9 downto 0);
    signal mulr_3_875 : std_logic_vector(9 downto 0);
    signal mulr_4_875 : std_logic_vector(9 downto 0);
    signal mulr_1_876 : std_logic_vector(9 downto 0);
    signal mulr_2_876 : std_logic_vector(9 downto 0);
    signal mulr_3_876 : std_logic_vector(9 downto 0);
    signal mulr_4_876 : std_logic_vector(9 downto 0);
    signal mulr_1_877 : std_logic_vector(9 downto 0);
    signal mulr_2_877 : std_logic_vector(9 downto 0);
    signal mulr_3_877 : std_logic_vector(9 downto 0);
    signal mulr_4_877 : std_logic_vector(9 downto 0);
    signal mulr_1_878 : std_logic_vector(9 downto 0);
    signal mulr_2_878 : std_logic_vector(9 downto 0);
    signal mulr_3_878 : std_logic_vector(9 downto 0);
    signal mulr_4_878 : std_logic_vector(9 downto 0);
    signal mulr_1_879 : std_logic_vector(9 downto 0);
    signal mulr_2_879 : std_logic_vector(9 downto 0);
    signal mulr_3_879 : std_logic_vector(9 downto 0);
    signal mulr_4_879 : std_logic_vector(9 downto 0);
    signal mulr_1_880 : std_logic_vector(9 downto 0);
    signal mulr_2_880 : std_logic_vector(9 downto 0);
    signal mulr_3_880 : std_logic_vector(9 downto 0);
    signal mulr_4_880 : std_logic_vector(9 downto 0);
    signal mulr_1_881 : std_logic_vector(9 downto 0);
    signal mulr_2_881 : std_logic_vector(9 downto 0);
    signal mulr_3_881 : std_logic_vector(9 downto 0);
    signal mulr_4_881 : std_logic_vector(9 downto 0);
    signal mulr_1_882 : std_logic_vector(9 downto 0);
    signal mulr_2_882 : std_logic_vector(9 downto 0);
    signal mulr_3_882 : std_logic_vector(9 downto 0);
    signal mulr_4_882 : std_logic_vector(9 downto 0);
    signal mulr_1_883 : std_logic_vector(9 downto 0);
    signal mulr_2_883 : std_logic_vector(9 downto 0);
    signal mulr_3_883 : std_logic_vector(9 downto 0);
    signal mulr_4_883 : std_logic_vector(9 downto 0);
    signal mulr_1_884 : std_logic_vector(9 downto 0);
    signal mulr_2_884 : std_logic_vector(9 downto 0);
    signal mulr_3_884 : std_logic_vector(9 downto 0);
    signal mulr_4_884 : std_logic_vector(9 downto 0);
    signal mulr_1_885 : std_logic_vector(9 downto 0);
    signal mulr_2_885 : std_logic_vector(9 downto 0);
    signal mulr_3_885 : std_logic_vector(9 downto 0);
    signal mulr_4_885 : std_logic_vector(9 downto 0);
    signal mulr_1_886 : std_logic_vector(9 downto 0);
    signal mulr_2_886 : std_logic_vector(9 downto 0);
    signal mulr_3_886 : std_logic_vector(9 downto 0);
    signal mulr_4_886 : std_logic_vector(9 downto 0);
    signal mulr_1_887 : std_logic_vector(9 downto 0);
    signal mulr_2_887 : std_logic_vector(9 downto 0);
    signal mulr_3_887 : std_logic_vector(9 downto 0);
    signal mulr_4_887 : std_logic_vector(9 downto 0);
    signal mulr_1_888 : std_logic_vector(9 downto 0);
    signal mulr_2_888 : std_logic_vector(9 downto 0);
    signal mulr_3_888 : std_logic_vector(9 downto 0);
    signal mulr_4_888 : std_logic_vector(9 downto 0);
    signal mulr_1_889 : std_logic_vector(9 downto 0);
    signal mulr_2_889 : std_logic_vector(9 downto 0);
    signal mulr_3_889 : std_logic_vector(9 downto 0);
    signal mulr_4_889 : std_logic_vector(9 downto 0);
    signal mulr_1_890 : std_logic_vector(9 downto 0);
    signal mulr_2_890 : std_logic_vector(9 downto 0);
    signal mulr_3_890 : std_logic_vector(9 downto 0);
    signal mulr_4_890 : std_logic_vector(9 downto 0);
    signal mulr_1_891 : std_logic_vector(9 downto 0);
    signal mulr_2_891 : std_logic_vector(9 downto 0);
    signal mulr_3_891 : std_logic_vector(9 downto 0);
    signal mulr_4_891 : std_logic_vector(9 downto 0);
    signal mulr_1_892 : std_logic_vector(9 downto 0);
    signal mulr_2_892 : std_logic_vector(9 downto 0);
    signal mulr_3_892 : std_logic_vector(9 downto 0);
    signal mulr_4_892 : std_logic_vector(9 downto 0);
    signal mulr_1_893 : std_logic_vector(9 downto 0);
    signal mulr_2_893 : std_logic_vector(9 downto 0);
    signal mulr_3_893 : std_logic_vector(9 downto 0);
    signal mulr_4_893 : std_logic_vector(9 downto 0);
    signal mulr_1_894 : std_logic_vector(9 downto 0);
    signal mulr_2_894 : std_logic_vector(9 downto 0);
    signal mulr_3_894 : std_logic_vector(9 downto 0);
    signal mulr_4_894 : std_logic_vector(9 downto 0);
    signal mulr_1_895 : std_logic_vector(9 downto 0);
    signal mulr_2_895 : std_logic_vector(9 downto 0);
    signal mulr_3_895 : std_logic_vector(9 downto 0);
    signal mulr_4_895 : std_logic_vector(9 downto 0);
    signal mulr_1_896 : std_logic_vector(9 downto 0);
    signal mulr_2_896 : std_logic_vector(9 downto 0);
    signal mulr_3_896 : std_logic_vector(9 downto 0);
    signal mulr_4_896 : std_logic_vector(9 downto 0);
    signal mulr_1_897 : std_logic_vector(9 downto 0);
    signal mulr_2_897 : std_logic_vector(9 downto 0);
    signal mulr_3_897 : std_logic_vector(9 downto 0);
    signal mulr_4_897 : std_logic_vector(9 downto 0);
    signal mulr_1_898 : std_logic_vector(9 downto 0);
    signal mulr_2_898 : std_logic_vector(9 downto 0);
    signal mulr_3_898 : std_logic_vector(9 downto 0);
    signal mulr_4_898 : std_logic_vector(9 downto 0);
    signal mulr_1_899 : std_logic_vector(9 downto 0);
    signal mulr_2_899 : std_logic_vector(9 downto 0);
    signal mulr_3_899 : std_logic_vector(9 downto 0);
    signal mulr_4_899 : std_logic_vector(9 downto 0);
    signal mulr_1_900 : std_logic_vector(9 downto 0);
    signal mulr_2_900 : std_logic_vector(9 downto 0);
    signal mulr_3_900 : std_logic_vector(9 downto 0);
    signal mulr_4_900 : std_logic_vector(9 downto 0);
    signal mulr_1_901 : std_logic_vector(9 downto 0);
    signal mulr_2_901 : std_logic_vector(9 downto 0);
    signal mulr_3_901 : std_logic_vector(9 downto 0);
    signal mulr_4_901 : std_logic_vector(9 downto 0);
    signal mulr_1_902 : std_logic_vector(9 downto 0);
    signal mulr_2_902 : std_logic_vector(9 downto 0);
    signal mulr_3_902 : std_logic_vector(9 downto 0);
    signal mulr_4_902 : std_logic_vector(9 downto 0);
    signal mulr_1_903 : std_logic_vector(9 downto 0);
    signal mulr_2_903 : std_logic_vector(9 downto 0);
    signal mulr_3_903 : std_logic_vector(9 downto 0);
    signal mulr_4_903 : std_logic_vector(9 downto 0);
    signal mulr_1_904 : std_logic_vector(9 downto 0);
    signal mulr_2_904 : std_logic_vector(9 downto 0);
    signal mulr_3_904 : std_logic_vector(9 downto 0);
    signal mulr_4_904 : std_logic_vector(9 downto 0);
    signal mulr_1_905 : std_logic_vector(9 downto 0);
    signal mulr_2_905 : std_logic_vector(9 downto 0);
    signal mulr_3_905 : std_logic_vector(9 downto 0);
    signal mulr_4_905 : std_logic_vector(9 downto 0);
    signal mulr_1_906 : std_logic_vector(9 downto 0);
    signal mulr_2_906 : std_logic_vector(9 downto 0);
    signal mulr_3_906 : std_logic_vector(9 downto 0);
    signal mulr_4_906 : std_logic_vector(9 downto 0);
    signal mulr_1_907 : std_logic_vector(9 downto 0);
    signal mulr_2_907 : std_logic_vector(9 downto 0);
    signal mulr_3_907 : std_logic_vector(9 downto 0);
    signal mulr_4_907 : std_logic_vector(9 downto 0);
    signal mulr_1_908 : std_logic_vector(9 downto 0);
    signal mulr_2_908 : std_logic_vector(9 downto 0);
    signal mulr_3_908 : std_logic_vector(9 downto 0);
    signal mulr_4_908 : std_logic_vector(9 downto 0);
    signal mulr_1_909 : std_logic_vector(9 downto 0);
    signal mulr_2_909 : std_logic_vector(9 downto 0);
    signal mulr_3_909 : std_logic_vector(9 downto 0);
    signal mulr_4_909 : std_logic_vector(9 downto 0);
    signal mulr_1_910 : std_logic_vector(9 downto 0);
    signal mulr_2_910 : std_logic_vector(9 downto 0);
    signal mulr_3_910 : std_logic_vector(9 downto 0);
    signal mulr_4_910 : std_logic_vector(9 downto 0);
    signal mulr_1_911 : std_logic_vector(9 downto 0);
    signal mulr_2_911 : std_logic_vector(9 downto 0);
    signal mulr_3_911 : std_logic_vector(9 downto 0);
    signal mulr_4_911 : std_logic_vector(9 downto 0);
    signal mulr_1_912 : std_logic_vector(9 downto 0);
    signal mulr_2_912 : std_logic_vector(9 downto 0);
    signal mulr_3_912 : std_logic_vector(9 downto 0);
    signal mulr_4_912 : std_logic_vector(9 downto 0);
    signal mulr_1_913 : std_logic_vector(9 downto 0);
    signal mulr_2_913 : std_logic_vector(9 downto 0);
    signal mulr_3_913 : std_logic_vector(9 downto 0);
    signal mulr_4_913 : std_logic_vector(9 downto 0);
    signal mulr_1_914 : std_logic_vector(9 downto 0);
    signal mulr_2_914 : std_logic_vector(9 downto 0);
    signal mulr_3_914 : std_logic_vector(9 downto 0);
    signal mulr_4_914 : std_logic_vector(9 downto 0);
    signal mulr_1_915 : std_logic_vector(9 downto 0);
    signal mulr_2_915 : std_logic_vector(9 downto 0);
    signal mulr_3_915 : std_logic_vector(9 downto 0);
    signal mulr_4_915 : std_logic_vector(9 downto 0);
    signal mulr_1_916 : std_logic_vector(9 downto 0);
    signal mulr_2_916 : std_logic_vector(9 downto 0);
    signal mulr_3_916 : std_logic_vector(9 downto 0);
    signal mulr_4_916 : std_logic_vector(9 downto 0);
    signal mulr_1_917 : std_logic_vector(9 downto 0);
    signal mulr_2_917 : std_logic_vector(9 downto 0);
    signal mulr_3_917 : std_logic_vector(9 downto 0);
    signal mulr_4_917 : std_logic_vector(9 downto 0);
    signal mulr_1_918 : std_logic_vector(9 downto 0);
    signal mulr_2_918 : std_logic_vector(9 downto 0);
    signal mulr_3_918 : std_logic_vector(9 downto 0);
    signal mulr_4_918 : std_logic_vector(9 downto 0);
    signal mulr_1_919 : std_logic_vector(9 downto 0);
    signal mulr_2_919 : std_logic_vector(9 downto 0);
    signal mulr_3_919 : std_logic_vector(9 downto 0);
    signal mulr_4_919 : std_logic_vector(9 downto 0);
    signal mulr_1_920 : std_logic_vector(9 downto 0);
    signal mulr_2_920 : std_logic_vector(9 downto 0);
    signal mulr_3_920 : std_logic_vector(9 downto 0);
    signal mulr_4_920 : std_logic_vector(9 downto 0);
    signal mulr_1_921 : std_logic_vector(9 downto 0);
    signal mulr_2_921 : std_logic_vector(9 downto 0);
    signal mulr_3_921 : std_logic_vector(9 downto 0);
    signal mulr_4_921 : std_logic_vector(9 downto 0);
    signal mulr_1_922 : std_logic_vector(9 downto 0);
    signal mulr_2_922 : std_logic_vector(9 downto 0);
    signal mulr_3_922 : std_logic_vector(9 downto 0);
    signal mulr_4_922 : std_logic_vector(9 downto 0);
    signal mulr_1_923 : std_logic_vector(9 downto 0);
    signal mulr_2_923 : std_logic_vector(9 downto 0);
    signal mulr_3_923 : std_logic_vector(9 downto 0);
    signal mulr_4_923 : std_logic_vector(9 downto 0);
    signal mulr_1_924 : std_logic_vector(9 downto 0);
    signal mulr_2_924 : std_logic_vector(9 downto 0);
    signal mulr_3_924 : std_logic_vector(9 downto 0);
    signal mulr_4_924 : std_logic_vector(9 downto 0);
    signal mulr_1_925 : std_logic_vector(9 downto 0);
    signal mulr_2_925 : std_logic_vector(9 downto 0);
    signal mulr_3_925 : std_logic_vector(9 downto 0);
    signal mulr_4_925 : std_logic_vector(9 downto 0);
    signal mulr_1_926 : std_logic_vector(9 downto 0);
    signal mulr_2_926 : std_logic_vector(9 downto 0);
    signal mulr_3_926 : std_logic_vector(9 downto 0);
    signal mulr_4_926 : std_logic_vector(9 downto 0);
    signal mulr_1_927 : std_logic_vector(9 downto 0);
    signal mulr_2_927 : std_logic_vector(9 downto 0);
    signal mulr_3_927 : std_logic_vector(9 downto 0);
    signal mulr_4_927 : std_logic_vector(9 downto 0);
    signal mulr_1_928 : std_logic_vector(9 downto 0);
    signal mulr_2_928 : std_logic_vector(9 downto 0);
    signal mulr_3_928 : std_logic_vector(9 downto 0);
    signal mulr_4_928 : std_logic_vector(9 downto 0);
    signal mulr_1_929 : std_logic_vector(9 downto 0);
    signal mulr_2_929 : std_logic_vector(9 downto 0);
    signal mulr_3_929 : std_logic_vector(9 downto 0);
    signal mulr_4_929 : std_logic_vector(9 downto 0);
    signal mulr_1_930 : std_logic_vector(9 downto 0);
    signal mulr_2_930 : std_logic_vector(9 downto 0);
    signal mulr_3_930 : std_logic_vector(9 downto 0);
    signal mulr_4_930 : std_logic_vector(9 downto 0);
    signal mulr_1_931 : std_logic_vector(9 downto 0);
    signal mulr_2_931 : std_logic_vector(9 downto 0);
    signal mulr_3_931 : std_logic_vector(9 downto 0);
    signal mulr_4_931 : std_logic_vector(9 downto 0);
    signal mulr_1_932 : std_logic_vector(9 downto 0);
    signal mulr_2_932 : std_logic_vector(9 downto 0);
    signal mulr_3_932 : std_logic_vector(9 downto 0);
    signal mulr_4_932 : std_logic_vector(9 downto 0);
    signal mulr_1_933 : std_logic_vector(9 downto 0);
    signal mulr_2_933 : std_logic_vector(9 downto 0);
    signal mulr_3_933 : std_logic_vector(9 downto 0);
    signal mulr_4_933 : std_logic_vector(9 downto 0);
    signal mulr_1_934 : std_logic_vector(9 downto 0);
    signal mulr_2_934 : std_logic_vector(9 downto 0);
    signal mulr_3_934 : std_logic_vector(9 downto 0);
    signal mulr_4_934 : std_logic_vector(9 downto 0);
    signal mulr_1_935 : std_logic_vector(9 downto 0);
    signal mulr_2_935 : std_logic_vector(9 downto 0);
    signal mulr_3_935 : std_logic_vector(9 downto 0);
    signal mulr_4_935 : std_logic_vector(9 downto 0);
    signal mulr_1_936 : std_logic_vector(9 downto 0);
    signal mulr_2_936 : std_logic_vector(9 downto 0);
    signal mulr_3_936 : std_logic_vector(9 downto 0);
    signal mulr_4_936 : std_logic_vector(9 downto 0);
    signal mulr_1_937 : std_logic_vector(9 downto 0);
    signal mulr_2_937 : std_logic_vector(9 downto 0);
    signal mulr_3_937 : std_logic_vector(9 downto 0);
    signal mulr_4_937 : std_logic_vector(9 downto 0);
    signal mulr_1_938 : std_logic_vector(9 downto 0);
    signal mulr_2_938 : std_logic_vector(9 downto 0);
    signal mulr_3_938 : std_logic_vector(9 downto 0);
    signal mulr_4_938 : std_logic_vector(9 downto 0);
    signal mulr_1_939 : std_logic_vector(9 downto 0);
    signal mulr_2_939 : std_logic_vector(9 downto 0);
    signal mulr_3_939 : std_logic_vector(9 downto 0);
    signal mulr_4_939 : std_logic_vector(9 downto 0);
    signal mulr_1_940 : std_logic_vector(9 downto 0);
    signal mulr_2_940 : std_logic_vector(9 downto 0);
    signal mulr_3_940 : std_logic_vector(9 downto 0);
    signal mulr_4_940 : std_logic_vector(9 downto 0);
    signal mulr_1_941 : std_logic_vector(9 downto 0);
    signal mulr_2_941 : std_logic_vector(9 downto 0);
    signal mulr_3_941 : std_logic_vector(9 downto 0);
    signal mulr_4_941 : std_logic_vector(9 downto 0);
    signal mulr_1_942 : std_logic_vector(9 downto 0);
    signal mulr_2_942 : std_logic_vector(9 downto 0);
    signal mulr_3_942 : std_logic_vector(9 downto 0);
    signal mulr_4_942 : std_logic_vector(9 downto 0);
    signal mulr_1_943 : std_logic_vector(9 downto 0);
    signal mulr_2_943 : std_logic_vector(9 downto 0);
    signal mulr_3_943 : std_logic_vector(9 downto 0);
    signal mulr_4_943 : std_logic_vector(9 downto 0);
    signal mulr_1_944 : std_logic_vector(9 downto 0);
    signal mulr_2_944 : std_logic_vector(9 downto 0);
    signal mulr_3_944 : std_logic_vector(9 downto 0);
    signal mulr_4_944 : std_logic_vector(9 downto 0);
    signal mulr_1_945 : std_logic_vector(9 downto 0);
    signal mulr_2_945 : std_logic_vector(9 downto 0);
    signal mulr_3_945 : std_logic_vector(9 downto 0);
    signal mulr_4_945 : std_logic_vector(9 downto 0);
    signal mulr_1_946 : std_logic_vector(9 downto 0);
    signal mulr_2_946 : std_logic_vector(9 downto 0);
    signal mulr_3_946 : std_logic_vector(9 downto 0);
    signal mulr_4_946 : std_logic_vector(9 downto 0);
    signal mulr_1_947 : std_logic_vector(9 downto 0);
    signal mulr_2_947 : std_logic_vector(9 downto 0);
    signal mulr_3_947 : std_logic_vector(9 downto 0);
    signal mulr_4_947 : std_logic_vector(9 downto 0);
    signal mulr_1_948 : std_logic_vector(9 downto 0);
    signal mulr_2_948 : std_logic_vector(9 downto 0);
    signal mulr_3_948 : std_logic_vector(9 downto 0);
    signal mulr_4_948 : std_logic_vector(9 downto 0);
    signal mulr_1_949 : std_logic_vector(9 downto 0);
    signal mulr_2_949 : std_logic_vector(9 downto 0);
    signal mulr_3_949 : std_logic_vector(9 downto 0);
    signal mulr_4_949 : std_logic_vector(9 downto 0);
    signal mulr_1_950 : std_logic_vector(9 downto 0);
    signal mulr_2_950 : std_logic_vector(9 downto 0);
    signal mulr_3_950 : std_logic_vector(9 downto 0);
    signal mulr_4_950 : std_logic_vector(9 downto 0);
    signal mulr_1_951 : std_logic_vector(9 downto 0);
    signal mulr_2_951 : std_logic_vector(9 downto 0);
    signal mulr_3_951 : std_logic_vector(9 downto 0);
    signal mulr_4_951 : std_logic_vector(9 downto 0);
    signal mulr_1_952 : std_logic_vector(9 downto 0);
    signal mulr_2_952 : std_logic_vector(9 downto 0);
    signal mulr_3_952 : std_logic_vector(9 downto 0);
    signal mulr_4_952 : std_logic_vector(9 downto 0);
    signal mulr_1_953 : std_logic_vector(9 downto 0);
    signal mulr_2_953 : std_logic_vector(9 downto 0);
    signal mulr_3_953 : std_logic_vector(9 downto 0);
    signal mulr_4_953 : std_logic_vector(9 downto 0);
    signal mulr_1_954 : std_logic_vector(9 downto 0);
    signal mulr_2_954 : std_logic_vector(9 downto 0);
    signal mulr_3_954 : std_logic_vector(9 downto 0);
    signal mulr_4_954 : std_logic_vector(9 downto 0);
    signal mulr_1_955 : std_logic_vector(9 downto 0);
    signal mulr_2_955 : std_logic_vector(9 downto 0);
    signal mulr_3_955 : std_logic_vector(9 downto 0);
    signal mulr_4_955 : std_logic_vector(9 downto 0);
    signal mulr_1_956 : std_logic_vector(9 downto 0);
    signal mulr_2_956 : std_logic_vector(9 downto 0);
    signal mulr_3_956 : std_logic_vector(9 downto 0);
    signal mulr_4_956 : std_logic_vector(9 downto 0);
    signal mulr_1_957 : std_logic_vector(9 downto 0);
    signal mulr_2_957 : std_logic_vector(9 downto 0);
    signal mulr_3_957 : std_logic_vector(9 downto 0);
    signal mulr_4_957 : std_logic_vector(9 downto 0);
    signal mulr_1_958 : std_logic_vector(9 downto 0);
    signal mulr_2_958 : std_logic_vector(9 downto 0);
    signal mulr_3_958 : std_logic_vector(9 downto 0);
    signal mulr_4_958 : std_logic_vector(9 downto 0);
    signal mulr_1_959 : std_logic_vector(9 downto 0);
    signal mulr_2_959 : std_logic_vector(9 downto 0);
    signal mulr_3_959 : std_logic_vector(9 downto 0);
    signal mulr_4_959 : std_logic_vector(9 downto 0);
    signal mulr_1_960 : std_logic_vector(9 downto 0);
    signal mulr_2_960 : std_logic_vector(9 downto 0);
    signal mulr_3_960 : std_logic_vector(9 downto 0);
    signal mulr_4_960 : std_logic_vector(9 downto 0);
    signal mulr_1_961 : std_logic_vector(9 downto 0);
    signal mulr_2_961 : std_logic_vector(9 downto 0);
    signal mulr_3_961 : std_logic_vector(9 downto 0);
    signal mulr_4_961 : std_logic_vector(9 downto 0);
    signal mulr_1_962 : std_logic_vector(9 downto 0);
    signal mulr_2_962 : std_logic_vector(9 downto 0);
    signal mulr_3_962 : std_logic_vector(9 downto 0);
    signal mulr_4_962 : std_logic_vector(9 downto 0);
    signal mulr_1_963 : std_logic_vector(9 downto 0);
    signal mulr_2_963 : std_logic_vector(9 downto 0);
    signal mulr_3_963 : std_logic_vector(9 downto 0);
    signal mulr_4_963 : std_logic_vector(9 downto 0);
    signal mulr_1_964 : std_logic_vector(9 downto 0);
    signal mulr_2_964 : std_logic_vector(9 downto 0);
    signal mulr_3_964 : std_logic_vector(9 downto 0);
    signal mulr_4_964 : std_logic_vector(9 downto 0);
    signal mulr_1_965 : std_logic_vector(9 downto 0);
    signal mulr_2_965 : std_logic_vector(9 downto 0);
    signal mulr_3_965 : std_logic_vector(9 downto 0);
    signal mulr_4_965 : std_logic_vector(9 downto 0);
    signal mulr_1_966 : std_logic_vector(9 downto 0);
    signal mulr_2_966 : std_logic_vector(9 downto 0);
    signal mulr_3_966 : std_logic_vector(9 downto 0);
    signal mulr_4_966 : std_logic_vector(9 downto 0);
    signal mulr_1_967 : std_logic_vector(9 downto 0);
    signal mulr_2_967 : std_logic_vector(9 downto 0);
    signal mulr_3_967 : std_logic_vector(9 downto 0);
    signal mulr_4_967 : std_logic_vector(9 downto 0);
    signal mulr_1_968 : std_logic_vector(9 downto 0);
    signal mulr_2_968 : std_logic_vector(9 downto 0);
    signal mulr_3_968 : std_logic_vector(9 downto 0);
    signal mulr_4_968 : std_logic_vector(9 downto 0);
    signal mulr_1_969 : std_logic_vector(9 downto 0);
    signal mulr_2_969 : std_logic_vector(9 downto 0);
    signal mulr_3_969 : std_logic_vector(9 downto 0);
    signal mulr_4_969 : std_logic_vector(9 downto 0);
    signal mulr_1_970 : std_logic_vector(9 downto 0);
    signal mulr_2_970 : std_logic_vector(9 downto 0);
    signal mulr_3_970 : std_logic_vector(9 downto 0);
    signal mulr_4_970 : std_logic_vector(9 downto 0);
    signal mulr_1_971 : std_logic_vector(9 downto 0);
    signal mulr_2_971 : std_logic_vector(9 downto 0);
    signal mulr_3_971 : std_logic_vector(9 downto 0);
    signal mulr_4_971 : std_logic_vector(9 downto 0);
    signal mulr_1_972 : std_logic_vector(9 downto 0);
    signal mulr_2_972 : std_logic_vector(9 downto 0);
    signal mulr_3_972 : std_logic_vector(9 downto 0);
    signal mulr_4_972 : std_logic_vector(9 downto 0);
    signal mulr_1_973 : std_logic_vector(9 downto 0);
    signal mulr_2_973 : std_logic_vector(9 downto 0);
    signal mulr_3_973 : std_logic_vector(9 downto 0);
    signal mulr_4_973 : std_logic_vector(9 downto 0);
    signal mulr_1_974 : std_logic_vector(9 downto 0);
    signal mulr_2_974 : std_logic_vector(9 downto 0);
    signal mulr_3_974 : std_logic_vector(9 downto 0);
    signal mulr_4_974 : std_logic_vector(9 downto 0);
    signal mulr_1_975 : std_logic_vector(9 downto 0);
    signal mulr_2_975 : std_logic_vector(9 downto 0);
    signal mulr_3_975 : std_logic_vector(9 downto 0);
    signal mulr_4_975 : std_logic_vector(9 downto 0);
    signal mulr_1_976 : std_logic_vector(9 downto 0);
    signal mulr_2_976 : std_logic_vector(9 downto 0);
    signal mulr_3_976 : std_logic_vector(9 downto 0);
    signal mulr_4_976 : std_logic_vector(9 downto 0);
    signal mulr_1_977 : std_logic_vector(9 downto 0);
    signal mulr_2_977 : std_logic_vector(9 downto 0);
    signal mulr_3_977 : std_logic_vector(9 downto 0);
    signal mulr_4_977 : std_logic_vector(9 downto 0);
    signal mulr_1_978 : std_logic_vector(9 downto 0);
    signal mulr_2_978 : std_logic_vector(9 downto 0);
    signal mulr_3_978 : std_logic_vector(9 downto 0);
    signal mulr_4_978 : std_logic_vector(9 downto 0);
    signal mulr_1_979 : std_logic_vector(9 downto 0);
    signal mulr_2_979 : std_logic_vector(9 downto 0);
    signal mulr_3_979 : std_logic_vector(9 downto 0);
    signal mulr_4_979 : std_logic_vector(9 downto 0);
    signal mulr_1_980 : std_logic_vector(9 downto 0);
    signal mulr_2_980 : std_logic_vector(9 downto 0);
    signal mulr_3_980 : std_logic_vector(9 downto 0);
    signal mulr_4_980 : std_logic_vector(9 downto 0);
    signal mulr_1_981 : std_logic_vector(9 downto 0);
    signal mulr_2_981 : std_logic_vector(9 downto 0);
    signal mulr_3_981 : std_logic_vector(9 downto 0);
    signal mulr_4_981 : std_logic_vector(9 downto 0);
    signal mulr_1_982 : std_logic_vector(9 downto 0);
    signal mulr_2_982 : std_logic_vector(9 downto 0);
    signal mulr_3_982 : std_logic_vector(9 downto 0);
    signal mulr_4_982 : std_logic_vector(9 downto 0);
    signal mulr_1_983 : std_logic_vector(9 downto 0);
    signal mulr_2_983 : std_logic_vector(9 downto 0);
    signal mulr_3_983 : std_logic_vector(9 downto 0);
    signal mulr_4_983 : std_logic_vector(9 downto 0);
    signal mulr_1_984 : std_logic_vector(9 downto 0);
    signal mulr_2_984 : std_logic_vector(9 downto 0);
    signal mulr_3_984 : std_logic_vector(9 downto 0);
    signal mulr_4_984 : std_logic_vector(9 downto 0);
    signal mulr_1_985 : std_logic_vector(9 downto 0);
    signal mulr_2_985 : std_logic_vector(9 downto 0);
    signal mulr_3_985 : std_logic_vector(9 downto 0);
    signal mulr_4_985 : std_logic_vector(9 downto 0);
    signal mulr_1_986 : std_logic_vector(9 downto 0);
    signal mulr_2_986 : std_logic_vector(9 downto 0);
    signal mulr_3_986 : std_logic_vector(9 downto 0);
    signal mulr_4_986 : std_logic_vector(9 downto 0);
    signal mulr_1_987 : std_logic_vector(9 downto 0);
    signal mulr_2_987 : std_logic_vector(9 downto 0);
    signal mulr_3_987 : std_logic_vector(9 downto 0);
    signal mulr_4_987 : std_logic_vector(9 downto 0);
    signal mulr_1_988 : std_logic_vector(9 downto 0);
    signal mulr_2_988 : std_logic_vector(9 downto 0);
    signal mulr_3_988 : std_logic_vector(9 downto 0);
    signal mulr_4_988 : std_logic_vector(9 downto 0);
    signal mulr_1_989 : std_logic_vector(9 downto 0);
    signal mulr_2_989 : std_logic_vector(9 downto 0);
    signal mulr_3_989 : std_logic_vector(9 downto 0);
    signal mulr_4_989 : std_logic_vector(9 downto 0);
    signal mulr_1_990 : std_logic_vector(9 downto 0);
    signal mulr_2_990 : std_logic_vector(9 downto 0);
    signal mulr_3_990 : std_logic_vector(9 downto 0);
    signal mulr_4_990 : std_logic_vector(9 downto 0);
    signal mulr_1_991 : std_logic_vector(9 downto 0);
    signal mulr_2_991 : std_logic_vector(9 downto 0);
    signal mulr_3_991 : std_logic_vector(9 downto 0);
    signal mulr_4_991 : std_logic_vector(9 downto 0);
    signal mulr_1_992 : std_logic_vector(9 downto 0);
    signal mulr_2_992 : std_logic_vector(9 downto 0);
    signal mulr_3_992 : std_logic_vector(9 downto 0);
    signal mulr_4_992 : std_logic_vector(9 downto 0);
    signal mulr_1_993 : std_logic_vector(9 downto 0);
    signal mulr_2_993 : std_logic_vector(9 downto 0);
    signal mulr_3_993 : std_logic_vector(9 downto 0);
    signal mulr_4_993 : std_logic_vector(9 downto 0);
    signal mulr_1_994 : std_logic_vector(9 downto 0);
    signal mulr_2_994 : std_logic_vector(9 downto 0);
    signal mulr_3_994 : std_logic_vector(9 downto 0);
    signal mulr_4_994 : std_logic_vector(9 downto 0);
    signal mulr_1_995 : std_logic_vector(9 downto 0);
    signal mulr_2_995 : std_logic_vector(9 downto 0);
    signal mulr_3_995 : std_logic_vector(9 downto 0);
    signal mulr_4_995 : std_logic_vector(9 downto 0);
    signal mulr_1_996 : std_logic_vector(9 downto 0);
    signal mulr_2_996 : std_logic_vector(9 downto 0);
    signal mulr_3_996 : std_logic_vector(9 downto 0);
    signal mulr_4_996 : std_logic_vector(9 downto 0);
    signal mulr_1_997 : std_logic_vector(9 downto 0);
    signal mulr_2_997 : std_logic_vector(9 downto 0);
    signal mulr_3_997 : std_logic_vector(9 downto 0);
    signal mulr_4_997 : std_logic_vector(9 downto 0);
    signal mulr_1_998 : std_logic_vector(9 downto 0);
    signal mulr_2_998 : std_logic_vector(9 downto 0);
    signal mulr_3_998 : std_logic_vector(9 downto 0);
    signal mulr_4_998 : std_logic_vector(9 downto 0);
    signal mulr_1_999 : std_logic_vector(9 downto 0);
    signal mulr_2_999 : std_logic_vector(9 downto 0);
    signal mulr_3_999 : std_logic_vector(9 downto 0);
    signal mulr_4_999 : std_logic_vector(9 downto 0);
    signal mulr_1_1000 : std_logic_vector(9 downto 0);
    signal mulr_2_1000 : std_logic_vector(9 downto 0);
    signal mulr_3_1000 : std_logic_vector(9 downto 0);
    signal mulr_4_1000 : std_logic_vector(9 downto 0);
    signal mulr_1_1001 : std_logic_vector(9 downto 0);
    signal mulr_2_1001 : std_logic_vector(9 downto 0);
    signal mulr_3_1001 : std_logic_vector(9 downto 0);
    signal mulr_4_1001 : std_logic_vector(9 downto 0);
    signal mulr_1_1002 : std_logic_vector(9 downto 0);
    signal mulr_2_1002 : std_logic_vector(9 downto 0);
    signal mulr_3_1002 : std_logic_vector(9 downto 0);
    signal mulr_4_1002 : std_logic_vector(9 downto 0);
    signal mulr_1_1003 : std_logic_vector(9 downto 0);
    signal mulr_2_1003 : std_logic_vector(9 downto 0);
    signal mulr_3_1003 : std_logic_vector(9 downto 0);
    signal mulr_4_1003 : std_logic_vector(9 downto 0);
    signal mulr_1_1004 : std_logic_vector(9 downto 0);
    signal mulr_2_1004 : std_logic_vector(9 downto 0);
    signal mulr_3_1004 : std_logic_vector(9 downto 0);
    signal mulr_4_1004 : std_logic_vector(9 downto 0);
    signal mulr_1_1005 : std_logic_vector(9 downto 0);
    signal mulr_2_1005 : std_logic_vector(9 downto 0);
    signal mulr_3_1005 : std_logic_vector(9 downto 0);
    signal mulr_4_1005 : std_logic_vector(9 downto 0);
    signal mulr_1_1006 : std_logic_vector(9 downto 0);
    signal mulr_2_1006 : std_logic_vector(9 downto 0);
    signal mulr_3_1006 : std_logic_vector(9 downto 0);
    signal mulr_4_1006 : std_logic_vector(9 downto 0);
    signal mulr_1_1007 : std_logic_vector(9 downto 0);
    signal mulr_2_1007 : std_logic_vector(9 downto 0);
    signal mulr_3_1007 : std_logic_vector(9 downto 0);
    signal mulr_4_1007 : std_logic_vector(9 downto 0);
    signal mulr_1_1008 : std_logic_vector(9 downto 0);
    signal mulr_2_1008 : std_logic_vector(9 downto 0);
    signal mulr_3_1008 : std_logic_vector(9 downto 0);
    signal mulr_4_1008 : std_logic_vector(9 downto 0);
    signal mulr_1_1009 : std_logic_vector(9 downto 0);
    signal mulr_2_1009 : std_logic_vector(9 downto 0);
    signal mulr_3_1009 : std_logic_vector(9 downto 0);
    signal mulr_4_1009 : std_logic_vector(9 downto 0);
    signal mulr_1_1010 : std_logic_vector(9 downto 0);
    signal mulr_2_1010 : std_logic_vector(9 downto 0);
    signal mulr_3_1010 : std_logic_vector(9 downto 0);
    signal mulr_4_1010 : std_logic_vector(9 downto 0);
    signal mulr_1_1011 : std_logic_vector(9 downto 0);
    signal mulr_2_1011 : std_logic_vector(9 downto 0);
    signal mulr_3_1011 : std_logic_vector(9 downto 0);
    signal mulr_4_1011 : std_logic_vector(9 downto 0);
    signal mulr_1_1012 : std_logic_vector(9 downto 0);
    signal mulr_2_1012 : std_logic_vector(9 downto 0);
    signal mulr_3_1012 : std_logic_vector(9 downto 0);
    signal mulr_4_1012 : std_logic_vector(9 downto 0);
    signal mulr_1_1013 : std_logic_vector(9 downto 0);
    signal mulr_2_1013 : std_logic_vector(9 downto 0);
    signal mulr_3_1013 : std_logic_vector(9 downto 0);
    signal mulr_4_1013 : std_logic_vector(9 downto 0);
    signal mulr_1_1014 : std_logic_vector(9 downto 0);
    signal mulr_2_1014 : std_logic_vector(9 downto 0);
    signal mulr_3_1014 : std_logic_vector(9 downto 0);
    signal mulr_4_1014 : std_logic_vector(9 downto 0);
    signal mulr_1_1015 : std_logic_vector(9 downto 0);
    signal mulr_2_1015 : std_logic_vector(9 downto 0);
    signal mulr_3_1015 : std_logic_vector(9 downto 0);
    signal mulr_4_1015 : std_logic_vector(9 downto 0);
    signal mulr_1_1016 : std_logic_vector(9 downto 0);
    signal mulr_2_1016 : std_logic_vector(9 downto 0);
    signal mulr_3_1016 : std_logic_vector(9 downto 0);
    signal mulr_4_1016 : std_logic_vector(9 downto 0);
    signal mulr_1_1017 : std_logic_vector(9 downto 0);
    signal mulr_2_1017 : std_logic_vector(9 downto 0);
    signal mulr_3_1017 : std_logic_vector(9 downto 0);
    signal mulr_4_1017 : std_logic_vector(9 downto 0);
    signal mulr_1_1018 : std_logic_vector(9 downto 0);
    signal mulr_2_1018 : std_logic_vector(9 downto 0);
    signal mulr_3_1018 : std_logic_vector(9 downto 0);
    signal mulr_4_1018 : std_logic_vector(9 downto 0);
    signal mulr_1_1019 : std_logic_vector(9 downto 0);
    signal mulr_2_1019 : std_logic_vector(9 downto 0);
    signal mulr_3_1019 : std_logic_vector(9 downto 0);
    signal mulr_4_1019 : std_logic_vector(9 downto 0);
    signal mulr_1_1020 : std_logic_vector(9 downto 0);
    signal mulr_2_1020 : std_logic_vector(9 downto 0);
    signal mulr_3_1020 : std_logic_vector(9 downto 0);
    signal mulr_4_1020 : std_logic_vector(9 downto 0);
    signal mulr_1_1021 : std_logic_vector(9 downto 0);
    signal mulr_2_1021 : std_logic_vector(9 downto 0);
    signal mulr_3_1021 : std_logic_vector(9 downto 0);
    signal mulr_4_1021 : std_logic_vector(9 downto 0);
    signal mulr_1_1022 : std_logic_vector(9 downto 0);
    signal mulr_2_1022 : std_logic_vector(9 downto 0);
    signal mulr_3_1022 : std_logic_vector(9 downto 0);
    signal mulr_4_1022 : std_logic_vector(9 downto 0);
    signal mulr_1_1023 : std_logic_vector(9 downto 0);
    signal mulr_2_1023 : std_logic_vector(9 downto 0);
    signal mulr_3_1023 : std_logic_vector(9 downto 0);
    signal mulr_4_1023 : std_logic_vector(9 downto 0);
    signal sumr_1 : std_logic_vector(9 downto 0);
    signal sumr_2 : std_logic_vector(9 downto 0);
    signal sumr_3 : std_logic_vector(9 downto 0);
    signal sumr_4 : std_logic_vector(9 downto 0);
    signal sumr_5 : std_logic_vector(9 downto 0);
    signal sumr_6 : std_logic_vector(9 downto 0);
    signal sumr_7 : std_logic_vector(9 downto 0);
    signal sumr_8 : std_logic_vector(9 downto 0);
    signal sumr_9 : std_logic_vector(9 downto 0);
    signal sumr_10 : std_logic_vector(9 downto 0);
    signal sumr_11 : std_logic_vector(9 downto 0);
    signal sumr_12 : std_logic_vector(9 downto 0);
    signal sumr_13 : std_logic_vector(9 downto 0);
    signal sumr_14 : std_logic_vector(9 downto 0);
    signal sumr_15 : std_logic_vector(9 downto 0);
    signal sumr_16 : std_logic_vector(9 downto 0);
    signal sumr_17 : std_logic_vector(9 downto 0);
    signal sumr_18 : std_logic_vector(9 downto 0);
    signal sumr_19 : std_logic_vector(9 downto 0);
    signal sumr_20 : std_logic_vector(9 downto 0);
    signal sumr_21 : std_logic_vector(9 downto 0);
    signal sumr_22 : std_logic_vector(9 downto 0);
    signal sumr_23 : std_logic_vector(9 downto 0);
    signal sumr_24 : std_logic_vector(9 downto 0);
    signal sumr_25 : std_logic_vector(9 downto 0);
    signal sumr_26 : std_logic_vector(9 downto 0);
    signal sumr_27 : std_logic_vector(9 downto 0);
    signal sumr_28 : std_logic_vector(9 downto 0);
    signal sumr_29 : std_logic_vector(9 downto 0);
    signal sumr_30 : std_logic_vector(9 downto 0);
    signal sumr_31 : std_logic_vector(9 downto 0);
    signal sumr_32 : std_logic_vector(9 downto 0);
    signal sumr_33 : std_logic_vector(9 downto 0);
    signal sumr_34 : std_logic_vector(9 downto 0);
    signal sumr_35 : std_logic_vector(9 downto 0);
    signal sumr_36 : std_logic_vector(9 downto 0);
    signal sumr_37 : std_logic_vector(9 downto 0);
    signal sumr_38 : std_logic_vector(9 downto 0);
    signal sumr_39 : std_logic_vector(9 downto 0);
    signal sumr_40 : std_logic_vector(9 downto 0);
    signal sumr_41 : std_logic_vector(9 downto 0);
    signal sumr_42 : std_logic_vector(9 downto 0);
    signal sumr_43 : std_logic_vector(9 downto 0);
    signal sumr_44 : std_logic_vector(9 downto 0);
    signal sumr_45 : std_logic_vector(9 downto 0);
    signal sumr_46 : std_logic_vector(9 downto 0);
    signal sumr_47 : std_logic_vector(9 downto 0);
    signal sumr_48 : std_logic_vector(9 downto 0);
    signal sumr_49 : std_logic_vector(9 downto 0);
    signal sumr_50 : std_logic_vector(9 downto 0);
    signal sumr_51 : std_logic_vector(9 downto 0);
    signal sumr_52 : std_logic_vector(9 downto 0);
    signal sumr_53 : std_logic_vector(9 downto 0);
    signal sumr_54 : std_logic_vector(9 downto 0);
    signal sumr_55 : std_logic_vector(9 downto 0);
    signal sumr_56 : std_logic_vector(9 downto 0);
    signal sumr_57 : std_logic_vector(9 downto 0);
    signal sumr_58 : std_logic_vector(9 downto 0);
    signal sumr_59 : std_logic_vector(9 downto 0);
    signal sumr_60 : std_logic_vector(9 downto 0);
    signal sumr_61 : std_logic_vector(9 downto 0);
    signal sumr_62 : std_logic_vector(9 downto 0);
    signal sumr_63 : std_logic_vector(9 downto 0);
    signal sumr_64 : std_logic_vector(9 downto 0);
    signal sumr_65 : std_logic_vector(9 downto 0);
    signal sumr_66 : std_logic_vector(9 downto 0);
    signal sumr_67 : std_logic_vector(9 downto 0);
    signal sumr_68 : std_logic_vector(9 downto 0);
    signal sumr_69 : std_logic_vector(9 downto 0);
    signal sumr_70 : std_logic_vector(9 downto 0);
    signal sumr_71 : std_logic_vector(9 downto 0);
    signal sumr_72 : std_logic_vector(9 downto 0);
    signal sumr_73 : std_logic_vector(9 downto 0);
    signal sumr_74 : std_logic_vector(9 downto 0);
    signal sumr_75 : std_logic_vector(9 downto 0);
    signal sumr_76 : std_logic_vector(9 downto 0);
    signal sumr_77 : std_logic_vector(9 downto 0);
    signal sumr_78 : std_logic_vector(9 downto 0);
    signal sumr_79 : std_logic_vector(9 downto 0);
    signal sumr_80 : std_logic_vector(9 downto 0);
    signal sumr_81 : std_logic_vector(9 downto 0);
    signal sumr_82 : std_logic_vector(9 downto 0);
    signal sumr_83 : std_logic_vector(9 downto 0);
    signal sumr_84 : std_logic_vector(9 downto 0);
    signal sumr_85 : std_logic_vector(9 downto 0);
    signal sumr_86 : std_logic_vector(9 downto 0);
    signal sumr_87 : std_logic_vector(9 downto 0);
    signal sumr_88 : std_logic_vector(9 downto 0);
    signal sumr_89 : std_logic_vector(9 downto 0);
    signal sumr_90 : std_logic_vector(9 downto 0);
    signal sumr_91 : std_logic_vector(9 downto 0);
    signal sumr_92 : std_logic_vector(9 downto 0);
    signal sumr_93 : std_logic_vector(9 downto 0);
    signal sumr_94 : std_logic_vector(9 downto 0);
    signal sumr_95 : std_logic_vector(9 downto 0);
    signal sumr_96 : std_logic_vector(9 downto 0);
    signal sumr_97 : std_logic_vector(9 downto 0);
    signal sumr_98 : std_logic_vector(9 downto 0);
    signal sumr_99 : std_logic_vector(9 downto 0);
    signal sumr_100 : std_logic_vector(9 downto 0);
    signal sumr_101 : std_logic_vector(9 downto 0);
    signal sumr_102 : std_logic_vector(9 downto 0);
    signal sumr_103 : std_logic_vector(9 downto 0);
    signal sumr_104 : std_logic_vector(9 downto 0);
    signal sumr_105 : std_logic_vector(9 downto 0);
    signal sumr_106 : std_logic_vector(9 downto 0);
    signal sumr_107 : std_logic_vector(9 downto 0);
    signal sumr_108 : std_logic_vector(9 downto 0);
    signal sumr_109 : std_logic_vector(9 downto 0);
    signal sumr_110 : std_logic_vector(9 downto 0);
    signal sumr_111 : std_logic_vector(9 downto 0);
    signal sumr_112 : std_logic_vector(9 downto 0);
    signal sumr_113 : std_logic_vector(9 downto 0);
    signal sumr_114 : std_logic_vector(9 downto 0);
    signal sumr_115 : std_logic_vector(9 downto 0);
    signal sumr_116 : std_logic_vector(9 downto 0);
    signal sumr_117 : std_logic_vector(9 downto 0);
    signal sumr_118 : std_logic_vector(9 downto 0);
    signal sumr_119 : std_logic_vector(9 downto 0);
    signal sumr_120 : std_logic_vector(9 downto 0);
    signal sumr_121 : std_logic_vector(9 downto 0);
    signal sumr_122 : std_logic_vector(9 downto 0);
    signal sumr_123 : std_logic_vector(9 downto 0);
    signal sumr_124 : std_logic_vector(9 downto 0);
    signal sumr_125 : std_logic_vector(9 downto 0);
    signal sumr_126 : std_logic_vector(9 downto 0);
    signal sumr_127 : std_logic_vector(9 downto 0);
    signal sumr_128 : std_logic_vector(9 downto 0);
    signal sumr_129 : std_logic_vector(9 downto 0);
    signal sumr_130 : std_logic_vector(9 downto 0);
    signal sumr_131 : std_logic_vector(9 downto 0);
    signal sumr_132 : std_logic_vector(9 downto 0);
    signal sumr_133 : std_logic_vector(9 downto 0);
    signal sumr_134 : std_logic_vector(9 downto 0);
    signal sumr_135 : std_logic_vector(9 downto 0);
    signal sumr_136 : std_logic_vector(9 downto 0);
    signal sumr_137 : std_logic_vector(9 downto 0);
    signal sumr_138 : std_logic_vector(9 downto 0);
    signal sumr_139 : std_logic_vector(9 downto 0);
    signal sumr_140 : std_logic_vector(9 downto 0);
    signal sumr_141 : std_logic_vector(9 downto 0);
    signal sumr_142 : std_logic_vector(9 downto 0);
    signal sumr_143 : std_logic_vector(9 downto 0);
    signal sumr_144 : std_logic_vector(9 downto 0);
    signal sumr_145 : std_logic_vector(9 downto 0);
    signal sumr_146 : std_logic_vector(9 downto 0);
    signal sumr_147 : std_logic_vector(9 downto 0);
    signal sumr_148 : std_logic_vector(9 downto 0);
    signal sumr_149 : std_logic_vector(9 downto 0);
    signal sumr_150 : std_logic_vector(9 downto 0);
    signal sumr_151 : std_logic_vector(9 downto 0);
    signal sumr_152 : std_logic_vector(9 downto 0);
    signal sumr_153 : std_logic_vector(9 downto 0);
    signal sumr_154 : std_logic_vector(9 downto 0);
    signal sumr_155 : std_logic_vector(9 downto 0);
    signal sumr_156 : std_logic_vector(9 downto 0);
    signal sumr_157 : std_logic_vector(9 downto 0);
    signal sumr_158 : std_logic_vector(9 downto 0);
    signal sumr_159 : std_logic_vector(9 downto 0);
    signal sumr_160 : std_logic_vector(9 downto 0);
    signal sumr_161 : std_logic_vector(9 downto 0);
    signal sumr_162 : std_logic_vector(9 downto 0);
    signal sumr_163 : std_logic_vector(9 downto 0);
    signal sumr_164 : std_logic_vector(9 downto 0);
    signal sumr_165 : std_logic_vector(9 downto 0);
    signal sumr_166 : std_logic_vector(9 downto 0);
    signal sumr_167 : std_logic_vector(9 downto 0);
    signal sumr_168 : std_logic_vector(9 downto 0);
    signal sumr_169 : std_logic_vector(9 downto 0);
    signal sumr_170 : std_logic_vector(9 downto 0);
    signal sumr_171 : std_logic_vector(9 downto 0);
    signal sumr_172 : std_logic_vector(9 downto 0);
    signal sumr_173 : std_logic_vector(9 downto 0);
    signal sumr_174 : std_logic_vector(9 downto 0);
    signal sumr_175 : std_logic_vector(9 downto 0);
    signal sumr_176 : std_logic_vector(9 downto 0);
    signal sumr_177 : std_logic_vector(9 downto 0);
    signal sumr_178 : std_logic_vector(9 downto 0);
    signal sumr_179 : std_logic_vector(9 downto 0);
    signal sumr_180 : std_logic_vector(9 downto 0);
    signal sumr_181 : std_logic_vector(9 downto 0);
    signal sumr_182 : std_logic_vector(9 downto 0);
    signal sumr_183 : std_logic_vector(9 downto 0);
    signal sumr_184 : std_logic_vector(9 downto 0);
    signal sumr_185 : std_logic_vector(9 downto 0);
    signal sumr_186 : std_logic_vector(9 downto 0);
    signal sumr_187 : std_logic_vector(9 downto 0);
    signal sumr_188 : std_logic_vector(9 downto 0);
    signal sumr_189 : std_logic_vector(9 downto 0);
    signal sumr_190 : std_logic_vector(9 downto 0);
    signal sumr_191 : std_logic_vector(9 downto 0);
    signal sumr_192 : std_logic_vector(9 downto 0);
    signal sumr_193 : std_logic_vector(9 downto 0);
    signal sumr_194 : std_logic_vector(9 downto 0);
    signal sumr_195 : std_logic_vector(9 downto 0);
    signal sumr_196 : std_logic_vector(9 downto 0);
    signal sumr_197 : std_logic_vector(9 downto 0);
    signal sumr_198 : std_logic_vector(9 downto 0);
    signal sumr_199 : std_logic_vector(9 downto 0);
    signal sumr_200 : std_logic_vector(9 downto 0);
    signal sumr_201 : std_logic_vector(9 downto 0);
    signal sumr_202 : std_logic_vector(9 downto 0);
    signal sumr_203 : std_logic_vector(9 downto 0);
    signal sumr_204 : std_logic_vector(9 downto 0);
    signal sumr_205 : std_logic_vector(9 downto 0);
    signal sumr_206 : std_logic_vector(9 downto 0);
    signal sumr_207 : std_logic_vector(9 downto 0);
    signal sumr_208 : std_logic_vector(9 downto 0);
    signal sumr_209 : std_logic_vector(9 downto 0);
    signal sumr_210 : std_logic_vector(9 downto 0);
    signal sumr_211 : std_logic_vector(9 downto 0);
    signal sumr_212 : std_logic_vector(9 downto 0);
    signal sumr_213 : std_logic_vector(9 downto 0);
    signal sumr_214 : std_logic_vector(9 downto 0);
    signal sumr_215 : std_logic_vector(9 downto 0);
    signal sumr_216 : std_logic_vector(9 downto 0);
    signal sumr_217 : std_logic_vector(9 downto 0);
    signal sumr_218 : std_logic_vector(9 downto 0);
    signal sumr_219 : std_logic_vector(9 downto 0);
    signal sumr_220 : std_logic_vector(9 downto 0);
    signal sumr_221 : std_logic_vector(9 downto 0);
    signal sumr_222 : std_logic_vector(9 downto 0);
    signal sumr_223 : std_logic_vector(9 downto 0);
    signal sumr_224 : std_logic_vector(9 downto 0);
    signal sumr_225 : std_logic_vector(9 downto 0);
    signal sumr_226 : std_logic_vector(9 downto 0);
    signal sumr_227 : std_logic_vector(9 downto 0);
    signal sumr_228 : std_logic_vector(9 downto 0);
    signal sumr_229 : std_logic_vector(9 downto 0);
    signal sumr_230 : std_logic_vector(9 downto 0);
    signal sumr_231 : std_logic_vector(9 downto 0);
    signal sumr_232 : std_logic_vector(9 downto 0);
    signal sumr_233 : std_logic_vector(9 downto 0);
    signal sumr_234 : std_logic_vector(9 downto 0);
    signal sumr_235 : std_logic_vector(9 downto 0);
    signal sumr_236 : std_logic_vector(9 downto 0);
    signal sumr_237 : std_logic_vector(9 downto 0);
    signal sumr_238 : std_logic_vector(9 downto 0);
    signal sumr_239 : std_logic_vector(9 downto 0);
    signal sumr_240 : std_logic_vector(9 downto 0);
    signal sumr_241 : std_logic_vector(9 downto 0);
    signal sumr_242 : std_logic_vector(9 downto 0);
    signal sumr_243 : std_logic_vector(9 downto 0);
    signal sumr_244 : std_logic_vector(9 downto 0);
    signal sumr_245 : std_logic_vector(9 downto 0);
    signal sumr_246 : std_logic_vector(9 downto 0);
    signal sumr_247 : std_logic_vector(9 downto 0);
    signal sumr_248 : std_logic_vector(9 downto 0);
    signal sumr_249 : std_logic_vector(9 downto 0);
    signal sumr_250 : std_logic_vector(9 downto 0);
    signal sumr_251 : std_logic_vector(9 downto 0);
    signal sumr_252 : std_logic_vector(9 downto 0);
    signal sumr_253 : std_logic_vector(9 downto 0);
    signal sumr_254 : std_logic_vector(9 downto 0);
    signal sumr_255 : std_logic_vector(9 downto 0);
    signal sumr_256 : std_logic_vector(9 downto 0);
    signal sumr_257 : std_logic_vector(9 downto 0);
    signal sumr_258 : std_logic_vector(9 downto 0);
    signal sumr_259 : std_logic_vector(9 downto 0);
    signal sumr_260 : std_logic_vector(9 downto 0);
    signal sumr_261 : std_logic_vector(9 downto 0);
    signal sumr_262 : std_logic_vector(9 downto 0);
    signal sumr_263 : std_logic_vector(9 downto 0);
    signal sumr_264 : std_logic_vector(9 downto 0);
    signal sumr_265 : std_logic_vector(9 downto 0);
    signal sumr_266 : std_logic_vector(9 downto 0);
    signal sumr_267 : std_logic_vector(9 downto 0);
    signal sumr_268 : std_logic_vector(9 downto 0);
    signal sumr_269 : std_logic_vector(9 downto 0);
    signal sumr_270 : std_logic_vector(9 downto 0);
    signal sumr_271 : std_logic_vector(9 downto 0);
    signal sumr_272 : std_logic_vector(9 downto 0);
    signal sumr_273 : std_logic_vector(9 downto 0);
    signal sumr_274 : std_logic_vector(9 downto 0);
    signal sumr_275 : std_logic_vector(9 downto 0);
    signal sumr_276 : std_logic_vector(9 downto 0);
    signal sumr_277 : std_logic_vector(9 downto 0);
    signal sumr_278 : std_logic_vector(9 downto 0);
    signal sumr_279 : std_logic_vector(9 downto 0);
    signal sumr_280 : std_logic_vector(9 downto 0);
    signal sumr_281 : std_logic_vector(9 downto 0);
    signal sumr_282 : std_logic_vector(9 downto 0);
    signal sumr_283 : std_logic_vector(9 downto 0);
    signal sumr_284 : std_logic_vector(9 downto 0);
    signal sumr_285 : std_logic_vector(9 downto 0);
    signal sumr_286 : std_logic_vector(9 downto 0);
    signal sumr_287 : std_logic_vector(9 downto 0);
    signal sumr_288 : std_logic_vector(9 downto 0);
    signal sumr_289 : std_logic_vector(9 downto 0);
    signal sumr_290 : std_logic_vector(9 downto 0);
    signal sumr_291 : std_logic_vector(9 downto 0);
    signal sumr_292 : std_logic_vector(9 downto 0);
    signal sumr_293 : std_logic_vector(9 downto 0);
    signal sumr_294 : std_logic_vector(9 downto 0);
    signal sumr_295 : std_logic_vector(9 downto 0);
    signal sumr_296 : std_logic_vector(9 downto 0);
    signal sumr_297 : std_logic_vector(9 downto 0);
    signal sumr_298 : std_logic_vector(9 downto 0);
    signal sumr_299 : std_logic_vector(9 downto 0);
    signal sumr_300 : std_logic_vector(9 downto 0);
    signal sumr_301 : std_logic_vector(9 downto 0);
    signal sumr_302 : std_logic_vector(9 downto 0);
    signal sumr_303 : std_logic_vector(9 downto 0);
    signal sumr_304 : std_logic_vector(9 downto 0);
    signal sumr_305 : std_logic_vector(9 downto 0);
    signal sumr_306 : std_logic_vector(9 downto 0);
    signal sumr_307 : std_logic_vector(9 downto 0);
    signal sumr_308 : std_logic_vector(9 downto 0);
    signal sumr_309 : std_logic_vector(9 downto 0);
    signal sumr_310 : std_logic_vector(9 downto 0);
    signal sumr_311 : std_logic_vector(9 downto 0);
    signal sumr_312 : std_logic_vector(9 downto 0);
    signal sumr_313 : std_logic_vector(9 downto 0);
    signal sumr_314 : std_logic_vector(9 downto 0);
    signal sumr_315 : std_logic_vector(9 downto 0);
    signal sumr_316 : std_logic_vector(9 downto 0);
    signal sumr_317 : std_logic_vector(9 downto 0);
    signal sumr_318 : std_logic_vector(9 downto 0);
    signal sumr_319 : std_logic_vector(9 downto 0);
    signal sumr_320 : std_logic_vector(9 downto 0);
    signal sumr_321 : std_logic_vector(9 downto 0);
    signal sumr_322 : std_logic_vector(9 downto 0);
    signal sumr_323 : std_logic_vector(9 downto 0);
    signal sumr_324 : std_logic_vector(9 downto 0);
    signal sumr_325 : std_logic_vector(9 downto 0);
    signal sumr_326 : std_logic_vector(9 downto 0);
    signal sumr_327 : std_logic_vector(9 downto 0);
    signal sumr_328 : std_logic_vector(9 downto 0);
    signal sumr_329 : std_logic_vector(9 downto 0);
    signal sumr_330 : std_logic_vector(9 downto 0);
    signal sumr_331 : std_logic_vector(9 downto 0);
    signal sumr_332 : std_logic_vector(9 downto 0);
    signal sumr_333 : std_logic_vector(9 downto 0);
    signal sumr_334 : std_logic_vector(9 downto 0);
    signal sumr_335 : std_logic_vector(9 downto 0);
    signal sumr_336 : std_logic_vector(9 downto 0);
    signal sumr_337 : std_logic_vector(9 downto 0);
    signal sumr_338 : std_logic_vector(9 downto 0);
    signal sumr_339 : std_logic_vector(9 downto 0);
    signal sumr_340 : std_logic_vector(9 downto 0);
    signal sumr_341 : std_logic_vector(9 downto 0);
    signal sumr_342 : std_logic_vector(9 downto 0);
    signal sumr_343 : std_logic_vector(9 downto 0);
    signal sumr_344 : std_logic_vector(9 downto 0);
    signal sumr_345 : std_logic_vector(9 downto 0);
    signal sumr_346 : std_logic_vector(9 downto 0);
    signal sumr_347 : std_logic_vector(9 downto 0);
    signal sumr_348 : std_logic_vector(9 downto 0);
    signal sumr_349 : std_logic_vector(9 downto 0);
    signal sumr_350 : std_logic_vector(9 downto 0);
    signal sumr_351 : std_logic_vector(9 downto 0);
    signal sumr_352 : std_logic_vector(9 downto 0);
    signal sumr_353 : std_logic_vector(9 downto 0);
    signal sumr_354 : std_logic_vector(9 downto 0);
    signal sumr_355 : std_logic_vector(9 downto 0);
    signal sumr_356 : std_logic_vector(9 downto 0);
    signal sumr_357 : std_logic_vector(9 downto 0);
    signal sumr_358 : std_logic_vector(9 downto 0);
    signal sumr_359 : std_logic_vector(9 downto 0);
    signal sumr_360 : std_logic_vector(9 downto 0);
    signal sumr_361 : std_logic_vector(9 downto 0);
    signal sumr_362 : std_logic_vector(9 downto 0);
    signal sumr_363 : std_logic_vector(9 downto 0);
    signal sumr_364 : std_logic_vector(9 downto 0);
    signal sumr_365 : std_logic_vector(9 downto 0);
    signal sumr_366 : std_logic_vector(9 downto 0);
    signal sumr_367 : std_logic_vector(9 downto 0);
    signal sumr_368 : std_logic_vector(9 downto 0);
    signal sumr_369 : std_logic_vector(9 downto 0);
    signal sumr_370 : std_logic_vector(9 downto 0);
    signal sumr_371 : std_logic_vector(9 downto 0);
    signal sumr_372 : std_logic_vector(9 downto 0);
    signal sumr_373 : std_logic_vector(9 downto 0);
    signal sumr_374 : std_logic_vector(9 downto 0);
    signal sumr_375 : std_logic_vector(9 downto 0);
    signal sumr_376 : std_logic_vector(9 downto 0);
    signal sumr_377 : std_logic_vector(9 downto 0);
    signal sumr_378 : std_logic_vector(9 downto 0);
    signal sumr_379 : std_logic_vector(9 downto 0);
    signal sumr_380 : std_logic_vector(9 downto 0);
    signal sumr_381 : std_logic_vector(9 downto 0);
    signal sumr_382 : std_logic_vector(9 downto 0);
    signal sumr_383 : std_logic_vector(9 downto 0);
    signal sumr_384 : std_logic_vector(9 downto 0);
    signal sumr_385 : std_logic_vector(9 downto 0);
    signal sumr_386 : std_logic_vector(9 downto 0);
    signal sumr_387 : std_logic_vector(9 downto 0);
    signal sumr_388 : std_logic_vector(9 downto 0);
    signal sumr_389 : std_logic_vector(9 downto 0);
    signal sumr_390 : std_logic_vector(9 downto 0);
    signal sumr_391 : std_logic_vector(9 downto 0);
    signal sumr_392 : std_logic_vector(9 downto 0);
    signal sumr_393 : std_logic_vector(9 downto 0);
    signal sumr_394 : std_logic_vector(9 downto 0);
    signal sumr_395 : std_logic_vector(9 downto 0);
    signal sumr_396 : std_logic_vector(9 downto 0);
    signal sumr_397 : std_logic_vector(9 downto 0);
    signal sumr_398 : std_logic_vector(9 downto 0);
    signal sumr_399 : std_logic_vector(9 downto 0);
    signal sumr_400 : std_logic_vector(9 downto 0);
    signal sumr_401 : std_logic_vector(9 downto 0);
    signal sumr_402 : std_logic_vector(9 downto 0);
    signal sumr_403 : std_logic_vector(9 downto 0);
    signal sumr_404 : std_logic_vector(9 downto 0);
    signal sumr_405 : std_logic_vector(9 downto 0);
    signal sumr_406 : std_logic_vector(9 downto 0);
    signal sumr_407 : std_logic_vector(9 downto 0);
    signal sumr_408 : std_logic_vector(9 downto 0);
    signal sumr_409 : std_logic_vector(9 downto 0);
    signal sumr_410 : std_logic_vector(9 downto 0);
    signal sumr_411 : std_logic_vector(9 downto 0);
    signal sumr_412 : std_logic_vector(9 downto 0);
    signal sumr_413 : std_logic_vector(9 downto 0);
    signal sumr_414 : std_logic_vector(9 downto 0);
    signal sumr_415 : std_logic_vector(9 downto 0);
    signal sumr_416 : std_logic_vector(9 downto 0);
    signal sumr_417 : std_logic_vector(9 downto 0);
    signal sumr_418 : std_logic_vector(9 downto 0);
    signal sumr_419 : std_logic_vector(9 downto 0);
    signal sumr_420 : std_logic_vector(9 downto 0);
    signal sumr_421 : std_logic_vector(9 downto 0);
    signal sumr_422 : std_logic_vector(9 downto 0);
    signal sumr_423 : std_logic_vector(9 downto 0);
    signal sumr_424 : std_logic_vector(9 downto 0);
    signal sumr_425 : std_logic_vector(9 downto 0);
    signal sumr_426 : std_logic_vector(9 downto 0);
    signal sumr_427 : std_logic_vector(9 downto 0);
    signal sumr_428 : std_logic_vector(9 downto 0);
    signal sumr_429 : std_logic_vector(9 downto 0);
    signal sumr_430 : std_logic_vector(9 downto 0);
    signal sumr_431 : std_logic_vector(9 downto 0);
    signal sumr_432 : std_logic_vector(9 downto 0);
    signal sumr_433 : std_logic_vector(9 downto 0);
    signal sumr_434 : std_logic_vector(9 downto 0);
    signal sumr_435 : std_logic_vector(9 downto 0);
    signal sumr_436 : std_logic_vector(9 downto 0);
    signal sumr_437 : std_logic_vector(9 downto 0);
    signal sumr_438 : std_logic_vector(9 downto 0);
    signal sumr_439 : std_logic_vector(9 downto 0);
    signal sumr_440 : std_logic_vector(9 downto 0);
    signal sumr_441 : std_logic_vector(9 downto 0);
    signal sumr_442 : std_logic_vector(9 downto 0);
    signal sumr_443 : std_logic_vector(9 downto 0);
    signal sumr_444 : std_logic_vector(9 downto 0);
    signal sumr_445 : std_logic_vector(9 downto 0);
    signal sumr_446 : std_logic_vector(9 downto 0);
    signal sumr_447 : std_logic_vector(9 downto 0);
    signal sumr_448 : std_logic_vector(9 downto 0);
    signal sumr_449 : std_logic_vector(9 downto 0);
    signal sumr_450 : std_logic_vector(9 downto 0);
    signal sumr_451 : std_logic_vector(9 downto 0);
    signal sumr_452 : std_logic_vector(9 downto 0);
    signal sumr_453 : std_logic_vector(9 downto 0);
    signal sumr_454 : std_logic_vector(9 downto 0);
    signal sumr_455 : std_logic_vector(9 downto 0);
    signal sumr_456 : std_logic_vector(9 downto 0);
    signal sumr_457 : std_logic_vector(9 downto 0);
    signal sumr_458 : std_logic_vector(9 downto 0);
    signal sumr_459 : std_logic_vector(9 downto 0);
    signal sumr_460 : std_logic_vector(9 downto 0);
    signal sumr_461 : std_logic_vector(9 downto 0);
    signal sumr_462 : std_logic_vector(9 downto 0);
    signal sumr_463 : std_logic_vector(9 downto 0);
    signal sumr_464 : std_logic_vector(9 downto 0);
    signal sumr_465 : std_logic_vector(9 downto 0);
    signal sumr_466 : std_logic_vector(9 downto 0);
    signal sumr_467 : std_logic_vector(9 downto 0);
    signal sumr_468 : std_logic_vector(9 downto 0);
    signal sumr_469 : std_logic_vector(9 downto 0);
    signal sumr_470 : std_logic_vector(9 downto 0);
    signal sumr_471 : std_logic_vector(9 downto 0);
    signal sumr_472 : std_logic_vector(9 downto 0);
    signal sumr_473 : std_logic_vector(9 downto 0);
    signal sumr_474 : std_logic_vector(9 downto 0);
    signal sumr_475 : std_logic_vector(9 downto 0);
    signal sumr_476 : std_logic_vector(9 downto 0);
    signal sumr_477 : std_logic_vector(9 downto 0);
    signal sumr_478 : std_logic_vector(9 downto 0);
    signal sumr_479 : std_logic_vector(9 downto 0);
    signal sumr_480 : std_logic_vector(9 downto 0);
    signal sumr_481 : std_logic_vector(9 downto 0);
    signal sumr_482 : std_logic_vector(9 downto 0);
    signal sumr_483 : std_logic_vector(9 downto 0);
    signal sumr_484 : std_logic_vector(9 downto 0);
    signal sumr_485 : std_logic_vector(9 downto 0);
    signal sumr_486 : std_logic_vector(9 downto 0);
    signal sumr_487 : std_logic_vector(9 downto 0);
    signal sumr_488 : std_logic_vector(9 downto 0);
    signal sumr_489 : std_logic_vector(9 downto 0);
    signal sumr_490 : std_logic_vector(9 downto 0);
    signal sumr_491 : std_logic_vector(9 downto 0);
    signal sumr_492 : std_logic_vector(9 downto 0);
    signal sumr_493 : std_logic_vector(9 downto 0);
    signal sumr_494 : std_logic_vector(9 downto 0);
    signal sumr_495 : std_logic_vector(9 downto 0);
    signal sumr_496 : std_logic_vector(9 downto 0);
    signal sumr_497 : std_logic_vector(9 downto 0);
    signal sumr_498 : std_logic_vector(9 downto 0);
    signal sumr_499 : std_logic_vector(9 downto 0);
    signal sumr_500 : std_logic_vector(9 downto 0);
    signal sumr_501 : std_logic_vector(9 downto 0);
    signal sumr_502 : std_logic_vector(9 downto 0);
    signal sumr_503 : std_logic_vector(9 downto 0);
    signal sumr_504 : std_logic_vector(9 downto 0);
    signal sumr_505 : std_logic_vector(9 downto 0);
    signal sumr_506 : std_logic_vector(9 downto 0);
    signal sumr_507 : std_logic_vector(9 downto 0);
    signal sumr_508 : std_logic_vector(9 downto 0);
    signal sumr_509 : std_logic_vector(9 downto 0);
    signal sumr_510 : std_logic_vector(9 downto 0);
    signal sumr_511 : std_logic_vector(9 downto 0);
    signal sumr_512 : std_logic_vector(9 downto 0);
    signal sumr_513 : std_logic_vector(9 downto 0);
    signal sumr_514 : std_logic_vector(9 downto 0);
    signal sumr_515 : std_logic_vector(9 downto 0);
    signal sumr_516 : std_logic_vector(9 downto 0);
    signal sumr_517 : std_logic_vector(9 downto 0);
    signal sumr_518 : std_logic_vector(9 downto 0);
    signal sumr_519 : std_logic_vector(9 downto 0);
    signal sumr_520 : std_logic_vector(9 downto 0);
    signal sumr_521 : std_logic_vector(9 downto 0);
    signal sumr_522 : std_logic_vector(9 downto 0);
    signal sumr_523 : std_logic_vector(9 downto 0);
    signal sumr_524 : std_logic_vector(9 downto 0);
    signal sumr_525 : std_logic_vector(9 downto 0);
    signal sumr_526 : std_logic_vector(9 downto 0);
    signal sumr_527 : std_logic_vector(9 downto 0);
    signal sumr_528 : std_logic_vector(9 downto 0);
    signal sumr_529 : std_logic_vector(9 downto 0);
    signal sumr_530 : std_logic_vector(9 downto 0);
    signal sumr_531 : std_logic_vector(9 downto 0);
    signal sumr_532 : std_logic_vector(9 downto 0);
    signal sumr_533 : std_logic_vector(9 downto 0);
    signal sumr_534 : std_logic_vector(9 downto 0);
    signal sumr_535 : std_logic_vector(9 downto 0);
    signal sumr_536 : std_logic_vector(9 downto 0);
    signal sumr_537 : std_logic_vector(9 downto 0);
    signal sumr_538 : std_logic_vector(9 downto 0);
    signal sumr_539 : std_logic_vector(9 downto 0);
    signal sumr_540 : std_logic_vector(9 downto 0);
    signal sumr_541 : std_logic_vector(9 downto 0);
    signal sumr_542 : std_logic_vector(9 downto 0);
    signal sumr_543 : std_logic_vector(9 downto 0);
    signal sumr_544 : std_logic_vector(9 downto 0);
    signal sumr_545 : std_logic_vector(9 downto 0);
    signal sumr_546 : std_logic_vector(9 downto 0);
    signal sumr_547 : std_logic_vector(9 downto 0);
    signal sumr_548 : std_logic_vector(9 downto 0);
    signal sumr_549 : std_logic_vector(9 downto 0);
    signal sumr_550 : std_logic_vector(9 downto 0);
    signal sumr_551 : std_logic_vector(9 downto 0);
    signal sumr_552 : std_logic_vector(9 downto 0);
    signal sumr_553 : std_logic_vector(9 downto 0);
    signal sumr_554 : std_logic_vector(9 downto 0);
    signal sumr_555 : std_logic_vector(9 downto 0);
    signal sumr_556 : std_logic_vector(9 downto 0);
    signal sumr_557 : std_logic_vector(9 downto 0);
    signal sumr_558 : std_logic_vector(9 downto 0);
    signal sumr_559 : std_logic_vector(9 downto 0);
    signal sumr_560 : std_logic_vector(9 downto 0);
    signal sumr_561 : std_logic_vector(9 downto 0);
    signal sumr_562 : std_logic_vector(9 downto 0);
    signal sumr_563 : std_logic_vector(9 downto 0);
    signal sumr_564 : std_logic_vector(9 downto 0);
    signal sumr_565 : std_logic_vector(9 downto 0);
    signal sumr_566 : std_logic_vector(9 downto 0);
    signal sumr_567 : std_logic_vector(9 downto 0);
    signal sumr_568 : std_logic_vector(9 downto 0);
    signal sumr_569 : std_logic_vector(9 downto 0);
    signal sumr_570 : std_logic_vector(9 downto 0);
    signal sumr_571 : std_logic_vector(9 downto 0);
    signal sumr_572 : std_logic_vector(9 downto 0);
    signal sumr_573 : std_logic_vector(9 downto 0);
    signal sumr_574 : std_logic_vector(9 downto 0);
    signal sumr_575 : std_logic_vector(9 downto 0);
    signal sumr_576 : std_logic_vector(9 downto 0);
    signal sumr_577 : std_logic_vector(9 downto 0);
    signal sumr_578 : std_logic_vector(9 downto 0);
    signal sumr_579 : std_logic_vector(9 downto 0);
    signal sumr_580 : std_logic_vector(9 downto 0);
    signal sumr_581 : std_logic_vector(9 downto 0);
    signal sumr_582 : std_logic_vector(9 downto 0);
    signal sumr_583 : std_logic_vector(9 downto 0);
    signal sumr_584 : std_logic_vector(9 downto 0);
    signal sumr_585 : std_logic_vector(9 downto 0);
    signal sumr_586 : std_logic_vector(9 downto 0);
    signal sumr_587 : std_logic_vector(9 downto 0);
    signal sumr_588 : std_logic_vector(9 downto 0);
    signal sumr_589 : std_logic_vector(9 downto 0);
    signal sumr_590 : std_logic_vector(9 downto 0);
    signal sumr_591 : std_logic_vector(9 downto 0);
    signal sumr_592 : std_logic_vector(9 downto 0);
    signal sumr_593 : std_logic_vector(9 downto 0);
    signal sumr_594 : std_logic_vector(9 downto 0);
    signal sumr_595 : std_logic_vector(9 downto 0);
    signal sumr_596 : std_logic_vector(9 downto 0);
    signal sumr_597 : std_logic_vector(9 downto 0);
    signal sumr_598 : std_logic_vector(9 downto 0);
    signal sumr_599 : std_logic_vector(9 downto 0);
    signal sumr_600 : std_logic_vector(9 downto 0);
    signal sumr_601 : std_logic_vector(9 downto 0);
    signal sumr_602 : std_logic_vector(9 downto 0);
    signal sumr_603 : std_logic_vector(9 downto 0);
    signal sumr_604 : std_logic_vector(9 downto 0);
    signal sumr_605 : std_logic_vector(9 downto 0);
    signal sumr_606 : std_logic_vector(9 downto 0);
    signal sumr_607 : std_logic_vector(9 downto 0);
    signal sumr_608 : std_logic_vector(9 downto 0);
    signal sumr_609 : std_logic_vector(9 downto 0);
    signal sumr_610 : std_logic_vector(9 downto 0);
    signal sumr_611 : std_logic_vector(9 downto 0);
    signal sumr_612 : std_logic_vector(9 downto 0);
    signal sumr_613 : std_logic_vector(9 downto 0);
    signal sumr_614 : std_logic_vector(9 downto 0);
    signal sumr_615 : std_logic_vector(9 downto 0);
    signal sumr_616 : std_logic_vector(9 downto 0);
    signal sumr_617 : std_logic_vector(9 downto 0);
    signal sumr_618 : std_logic_vector(9 downto 0);
    signal sumr_619 : std_logic_vector(9 downto 0);
    signal sumr_620 : std_logic_vector(9 downto 0);
    signal sumr_621 : std_logic_vector(9 downto 0);
    signal sumr_622 : std_logic_vector(9 downto 0);
    signal sumr_623 : std_logic_vector(9 downto 0);
    signal sumr_624 : std_logic_vector(9 downto 0);
    signal sumr_625 : std_logic_vector(9 downto 0);
    signal sumr_626 : std_logic_vector(9 downto 0);
    signal sumr_627 : std_logic_vector(9 downto 0);
    signal sumr_628 : std_logic_vector(9 downto 0);
    signal sumr_629 : std_logic_vector(9 downto 0);
    signal sumr_630 : std_logic_vector(9 downto 0);
    signal sumr_631 : std_logic_vector(9 downto 0);
    signal sumr_632 : std_logic_vector(9 downto 0);
    signal sumr_633 : std_logic_vector(9 downto 0);
    signal sumr_634 : std_logic_vector(9 downto 0);
    signal sumr_635 : std_logic_vector(9 downto 0);
    signal sumr_636 : std_logic_vector(9 downto 0);
    signal sumr_637 : std_logic_vector(9 downto 0);
    signal sumr_638 : std_logic_vector(9 downto 0);
    signal sumr_639 : std_logic_vector(9 downto 0);
    signal sumr_640 : std_logic_vector(9 downto 0);
    signal sumr_641 : std_logic_vector(9 downto 0);
    signal sumr_642 : std_logic_vector(9 downto 0);
    signal sumr_643 : std_logic_vector(9 downto 0);
    signal sumr_644 : std_logic_vector(9 downto 0);
    signal sumr_645 : std_logic_vector(9 downto 0);
    signal sumr_646 : std_logic_vector(9 downto 0);
    signal sumr_647 : std_logic_vector(9 downto 0);
    signal sumr_648 : std_logic_vector(9 downto 0);
    signal sumr_649 : std_logic_vector(9 downto 0);
    signal sumr_650 : std_logic_vector(9 downto 0);
    signal sumr_651 : std_logic_vector(9 downto 0);
    signal sumr_652 : std_logic_vector(9 downto 0);
    signal sumr_653 : std_logic_vector(9 downto 0);
    signal sumr_654 : std_logic_vector(9 downto 0);
    signal sumr_655 : std_logic_vector(9 downto 0);
    signal sumr_656 : std_logic_vector(9 downto 0);
    signal sumr_657 : std_logic_vector(9 downto 0);
    signal sumr_658 : std_logic_vector(9 downto 0);
    signal sumr_659 : std_logic_vector(9 downto 0);
    signal sumr_660 : std_logic_vector(9 downto 0);
    signal sumr_661 : std_logic_vector(9 downto 0);
    signal sumr_662 : std_logic_vector(9 downto 0);
    signal sumr_663 : std_logic_vector(9 downto 0);
    signal sumr_664 : std_logic_vector(9 downto 0);
    signal sumr_665 : std_logic_vector(9 downto 0);
    signal sumr_666 : std_logic_vector(9 downto 0);
    signal sumr_667 : std_logic_vector(9 downto 0);
    signal sumr_668 : std_logic_vector(9 downto 0);
    signal sumr_669 : std_logic_vector(9 downto 0);
    signal sumr_670 : std_logic_vector(9 downto 0);
    signal sumr_671 : std_logic_vector(9 downto 0);
    signal sumr_672 : std_logic_vector(9 downto 0);
    signal sumr_673 : std_logic_vector(9 downto 0);
    signal sumr_674 : std_logic_vector(9 downto 0);
    signal sumr_675 : std_logic_vector(9 downto 0);
    signal sumr_676 : std_logic_vector(9 downto 0);
    signal sumr_677 : std_logic_vector(9 downto 0);
    signal sumr_678 : std_logic_vector(9 downto 0);
    signal sumr_679 : std_logic_vector(9 downto 0);
    signal sumr_680 : std_logic_vector(9 downto 0);
    signal sumr_681 : std_logic_vector(9 downto 0);
    signal sumr_682 : std_logic_vector(9 downto 0);
    signal sumr_683 : std_logic_vector(9 downto 0);
    signal sumr_684 : std_logic_vector(9 downto 0);
    signal sumr_685 : std_logic_vector(9 downto 0);
    signal sumr_686 : std_logic_vector(9 downto 0);
    signal sumr_687 : std_logic_vector(9 downto 0);
    signal sumr_688 : std_logic_vector(9 downto 0);
    signal sumr_689 : std_logic_vector(9 downto 0);
    signal sumr_690 : std_logic_vector(9 downto 0);
    signal sumr_691 : std_logic_vector(9 downto 0);
    signal sumr_692 : std_logic_vector(9 downto 0);
    signal sumr_693 : std_logic_vector(9 downto 0);
    signal sumr_694 : std_logic_vector(9 downto 0);
    signal sumr_695 : std_logic_vector(9 downto 0);
    signal sumr_696 : std_logic_vector(9 downto 0);
    signal sumr_697 : std_logic_vector(9 downto 0);
    signal sumr_698 : std_logic_vector(9 downto 0);
    signal sumr_699 : std_logic_vector(9 downto 0);
    signal sumr_700 : std_logic_vector(9 downto 0);
    signal sumr_701 : std_logic_vector(9 downto 0);
    signal sumr_702 : std_logic_vector(9 downto 0);
    signal sumr_703 : std_logic_vector(9 downto 0);
    signal sumr_704 : std_logic_vector(9 downto 0);
    signal sumr_705 : std_logic_vector(9 downto 0);
    signal sumr_706 : std_logic_vector(9 downto 0);
    signal sumr_707 : std_logic_vector(9 downto 0);
    signal sumr_708 : std_logic_vector(9 downto 0);
    signal sumr_709 : std_logic_vector(9 downto 0);
    signal sumr_710 : std_logic_vector(9 downto 0);
    signal sumr_711 : std_logic_vector(9 downto 0);
    signal sumr_712 : std_logic_vector(9 downto 0);
    signal sumr_713 : std_logic_vector(9 downto 0);
    signal sumr_714 : std_logic_vector(9 downto 0);
    signal sumr_715 : std_logic_vector(9 downto 0);
    signal sumr_716 : std_logic_vector(9 downto 0);
    signal sumr_717 : std_logic_vector(9 downto 0);
    signal sumr_718 : std_logic_vector(9 downto 0);
    signal sumr_719 : std_logic_vector(9 downto 0);
    signal sumr_720 : std_logic_vector(9 downto 0);
    signal sumr_721 : std_logic_vector(9 downto 0);
    signal sumr_722 : std_logic_vector(9 downto 0);
    signal sumr_723 : std_logic_vector(9 downto 0);
    signal sumr_724 : std_logic_vector(9 downto 0);
    signal sumr_725 : std_logic_vector(9 downto 0);
    signal sumr_726 : std_logic_vector(9 downto 0);
    signal sumr_727 : std_logic_vector(9 downto 0);
    signal sumr_728 : std_logic_vector(9 downto 0);
    signal sumr_729 : std_logic_vector(9 downto 0);
    signal sumr_730 : std_logic_vector(9 downto 0);
    signal sumr_731 : std_logic_vector(9 downto 0);
    signal sumr_732 : std_logic_vector(9 downto 0);
    signal sumr_733 : std_logic_vector(9 downto 0);
    signal sumr_734 : std_logic_vector(9 downto 0);
    signal sumr_735 : std_logic_vector(9 downto 0);
    signal sumr_736 : std_logic_vector(9 downto 0);
    signal sumr_737 : std_logic_vector(9 downto 0);
    signal sumr_738 : std_logic_vector(9 downto 0);
    signal sumr_739 : std_logic_vector(9 downto 0);
    signal sumr_740 : std_logic_vector(9 downto 0);
    signal sumr_741 : std_logic_vector(9 downto 0);
    signal sumr_742 : std_logic_vector(9 downto 0);
    signal sumr_743 : std_logic_vector(9 downto 0);
    signal sumr_744 : std_logic_vector(9 downto 0);
    signal sumr_745 : std_logic_vector(9 downto 0);
    signal sumr_746 : std_logic_vector(9 downto 0);
    signal sumr_747 : std_logic_vector(9 downto 0);
    signal sumr_748 : std_logic_vector(9 downto 0);
    signal sumr_749 : std_logic_vector(9 downto 0);
    signal sumr_750 : std_logic_vector(9 downto 0);
    signal sumr_751 : std_logic_vector(9 downto 0);
    signal sumr_752 : std_logic_vector(9 downto 0);
    signal sumr_753 : std_logic_vector(9 downto 0);
    signal sumr_754 : std_logic_vector(9 downto 0);
    signal sumr_755 : std_logic_vector(9 downto 0);
    signal sumr_756 : std_logic_vector(9 downto 0);
    signal sumr_757 : std_logic_vector(9 downto 0);
    signal sumr_758 : std_logic_vector(9 downto 0);
    signal sumr_759 : std_logic_vector(9 downto 0);
    signal sumr_760 : std_logic_vector(9 downto 0);
    signal sumr_761 : std_logic_vector(9 downto 0);
    signal sumr_762 : std_logic_vector(9 downto 0);
    signal sumr_763 : std_logic_vector(9 downto 0);
    signal sumr_764 : std_logic_vector(9 downto 0);
    signal sumr_765 : std_logic_vector(9 downto 0);
    signal sumr_766 : std_logic_vector(9 downto 0);
    signal sumr_767 : std_logic_vector(9 downto 0);
    signal sumr_768 : std_logic_vector(9 downto 0);
    signal sumr_769 : std_logic_vector(9 downto 0);
    signal sumr_770 : std_logic_vector(9 downto 0);
    signal sumr_771 : std_logic_vector(9 downto 0);
    signal sumr_772 : std_logic_vector(9 downto 0);
    signal sumr_773 : std_logic_vector(9 downto 0);
    signal sumr_774 : std_logic_vector(9 downto 0);
    signal sumr_775 : std_logic_vector(9 downto 0);
    signal sumr_776 : std_logic_vector(9 downto 0);
    signal sumr_777 : std_logic_vector(9 downto 0);
    signal sumr_778 : std_logic_vector(9 downto 0);
    signal sumr_779 : std_logic_vector(9 downto 0);
    signal sumr_780 : std_logic_vector(9 downto 0);
    signal sumr_781 : std_logic_vector(9 downto 0);
    signal sumr_782 : std_logic_vector(9 downto 0);
    signal sumr_783 : std_logic_vector(9 downto 0);
    signal sumr_784 : std_logic_vector(9 downto 0);
    signal sumr_785 : std_logic_vector(9 downto 0);
    signal sumr_786 : std_logic_vector(9 downto 0);
    signal sumr_787 : std_logic_vector(9 downto 0);
    signal sumr_788 : std_logic_vector(9 downto 0);
    signal sumr_789 : std_logic_vector(9 downto 0);
    signal sumr_790 : std_logic_vector(9 downto 0);
    signal sumr_791 : std_logic_vector(9 downto 0);
    signal sumr_792 : std_logic_vector(9 downto 0);
    signal sumr_793 : std_logic_vector(9 downto 0);
    signal sumr_794 : std_logic_vector(9 downto 0);
    signal sumr_795 : std_logic_vector(9 downto 0);
    signal sumr_796 : std_logic_vector(9 downto 0);
    signal sumr_797 : std_logic_vector(9 downto 0);
    signal sumr_798 : std_logic_vector(9 downto 0);
    signal sumr_799 : std_logic_vector(9 downto 0);
    signal sumr_800 : std_logic_vector(9 downto 0);
    signal sumr_801 : std_logic_vector(9 downto 0);
    signal sumr_802 : std_logic_vector(9 downto 0);
    signal sumr_803 : std_logic_vector(9 downto 0);
    signal sumr_804 : std_logic_vector(9 downto 0);
    signal sumr_805 : std_logic_vector(9 downto 0);
    signal sumr_806 : std_logic_vector(9 downto 0);
    signal sumr_807 : std_logic_vector(9 downto 0);
    signal sumr_808 : std_logic_vector(9 downto 0);
    signal sumr_809 : std_logic_vector(9 downto 0);
    signal sumr_810 : std_logic_vector(9 downto 0);
    signal sumr_811 : std_logic_vector(9 downto 0);
    signal sumr_812 : std_logic_vector(9 downto 0);
    signal sumr_813 : std_logic_vector(9 downto 0);
    signal sumr_814 : std_logic_vector(9 downto 0);
    signal sumr_815 : std_logic_vector(9 downto 0);
    signal sumr_816 : std_logic_vector(9 downto 0);
    signal sumr_817 : std_logic_vector(9 downto 0);
    signal sumr_818 : std_logic_vector(9 downto 0);
    signal sumr_819 : std_logic_vector(9 downto 0);
    signal sumr_820 : std_logic_vector(9 downto 0);
    signal sumr_821 : std_logic_vector(9 downto 0);
    signal sumr_822 : std_logic_vector(9 downto 0);
    signal sumr_823 : std_logic_vector(9 downto 0);
    signal sumr_824 : std_logic_vector(9 downto 0);
    signal sumr_825 : std_logic_vector(9 downto 0);
    signal sumr_826 : std_logic_vector(9 downto 0);
    signal sumr_827 : std_logic_vector(9 downto 0);
    signal sumr_828 : std_logic_vector(9 downto 0);
    signal sumr_829 : std_logic_vector(9 downto 0);
    signal sumr_830 : std_logic_vector(9 downto 0);
    signal sumr_831 : std_logic_vector(9 downto 0);
    signal sumr_832 : std_logic_vector(9 downto 0);
    signal sumr_833 : std_logic_vector(9 downto 0);
    signal sumr_834 : std_logic_vector(9 downto 0);
    signal sumr_835 : std_logic_vector(9 downto 0);
    signal sumr_836 : std_logic_vector(9 downto 0);
    signal sumr_837 : std_logic_vector(9 downto 0);
    signal sumr_838 : std_logic_vector(9 downto 0);
    signal sumr_839 : std_logic_vector(9 downto 0);
    signal sumr_840 : std_logic_vector(9 downto 0);
    signal sumr_841 : std_logic_vector(9 downto 0);
    signal sumr_842 : std_logic_vector(9 downto 0);
    signal sumr_843 : std_logic_vector(9 downto 0);
    signal sumr_844 : std_logic_vector(9 downto 0);
    signal sumr_845 : std_logic_vector(9 downto 0);
    signal sumr_846 : std_logic_vector(9 downto 0);
    signal sumr_847 : std_logic_vector(9 downto 0);
    signal sumr_848 : std_logic_vector(9 downto 0);
    signal sumr_849 : std_logic_vector(9 downto 0);
    signal sumr_850 : std_logic_vector(9 downto 0);
    signal sumr_851 : std_logic_vector(9 downto 0);
    signal sumr_852 : std_logic_vector(9 downto 0);
    signal sumr_853 : std_logic_vector(9 downto 0);
    signal sumr_854 : std_logic_vector(9 downto 0);
    signal sumr_855 : std_logic_vector(9 downto 0);
    signal sumr_856 : std_logic_vector(9 downto 0);
    signal sumr_857 : std_logic_vector(9 downto 0);
    signal sumr_858 : std_logic_vector(9 downto 0);
    signal sumr_859 : std_logic_vector(9 downto 0);
    signal sumr_860 : std_logic_vector(9 downto 0);
    signal sumr_861 : std_logic_vector(9 downto 0);
    signal sumr_862 : std_logic_vector(9 downto 0);
    signal sumr_863 : std_logic_vector(9 downto 0);
    signal sumr_864 : std_logic_vector(9 downto 0);
    signal sumr_865 : std_logic_vector(9 downto 0);
    signal sumr_866 : std_logic_vector(9 downto 0);
    signal sumr_867 : std_logic_vector(9 downto 0);
    signal sumr_868 : std_logic_vector(9 downto 0);
    signal sumr_869 : std_logic_vector(9 downto 0);
    signal sumr_870 : std_logic_vector(9 downto 0);
    signal sumr_871 : std_logic_vector(9 downto 0);
    signal sumr_872 : std_logic_vector(9 downto 0);
    signal sumr_873 : std_logic_vector(9 downto 0);
    signal sumr_874 : std_logic_vector(9 downto 0);
    signal sumr_875 : std_logic_vector(9 downto 0);
    signal sumr_876 : std_logic_vector(9 downto 0);
    signal sumr_877 : std_logic_vector(9 downto 0);
    signal sumr_878 : std_logic_vector(9 downto 0);
    signal sumr_879 : std_logic_vector(9 downto 0);
    signal sumr_880 : std_logic_vector(9 downto 0);
    signal sumr_881 : std_logic_vector(9 downto 0);
    signal sumr_882 : std_logic_vector(9 downto 0);
    signal sumr_883 : std_logic_vector(9 downto 0);
    signal sumr_884 : std_logic_vector(9 downto 0);
    signal sumr_885 : std_logic_vector(9 downto 0);
    signal sumr_886 : std_logic_vector(9 downto 0);
    signal sumr_887 : std_logic_vector(9 downto 0);
    signal sumr_888 : std_logic_vector(9 downto 0);
    signal sumr_889 : std_logic_vector(9 downto 0);
    signal sumr_890 : std_logic_vector(9 downto 0);
    signal sumr_891 : std_logic_vector(9 downto 0);
    signal sumr_892 : std_logic_vector(9 downto 0);
    signal sumr_893 : std_logic_vector(9 downto 0);
    signal sumr_894 : std_logic_vector(9 downto 0);
    signal sumr_895 : std_logic_vector(9 downto 0);
    signal sumr_896 : std_logic_vector(9 downto 0);
    signal sumr_897 : std_logic_vector(9 downto 0);
    signal sumr_898 : std_logic_vector(9 downto 0);
    signal sumr_899 : std_logic_vector(9 downto 0);
    signal sumr_900 : std_logic_vector(9 downto 0);
    signal sumr_901 : std_logic_vector(9 downto 0);
    signal sumr_902 : std_logic_vector(9 downto 0);
    signal sumr_903 : std_logic_vector(9 downto 0);
    signal sumr_904 : std_logic_vector(9 downto 0);
    signal sumr_905 : std_logic_vector(9 downto 0);
    signal sumr_906 : std_logic_vector(9 downto 0);
    signal sumr_907 : std_logic_vector(9 downto 0);
    signal sumr_908 : std_logic_vector(9 downto 0);
    signal sumr_909 : std_logic_vector(9 downto 0);
    signal sumr_910 : std_logic_vector(9 downto 0);
    signal sumr_911 : std_logic_vector(9 downto 0);
    signal sumr_912 : std_logic_vector(9 downto 0);
    signal sumr_913 : std_logic_vector(9 downto 0);
    signal sumr_914 : std_logic_vector(9 downto 0);
    signal sumr_915 : std_logic_vector(9 downto 0);
    signal sumr_916 : std_logic_vector(9 downto 0);
    signal sumr_917 : std_logic_vector(9 downto 0);
    signal sumr_918 : std_logic_vector(9 downto 0);
    signal sumr_919 : std_logic_vector(9 downto 0);
    signal sumr_920 : std_logic_vector(9 downto 0);
    signal sumr_921 : std_logic_vector(9 downto 0);
    signal sumr_922 : std_logic_vector(9 downto 0);
    signal sumr_923 : std_logic_vector(9 downto 0);
    signal sumr_924 : std_logic_vector(9 downto 0);
    signal sumr_925 : std_logic_vector(9 downto 0);
    signal sumr_926 : std_logic_vector(9 downto 0);
    signal sumr_927 : std_logic_vector(9 downto 0);
    signal sumr_928 : std_logic_vector(9 downto 0);
    signal sumr_929 : std_logic_vector(9 downto 0);
    signal sumr_930 : std_logic_vector(9 downto 0);
    signal sumr_931 : std_logic_vector(9 downto 0);
    signal sumr_932 : std_logic_vector(9 downto 0);
    signal sumr_933 : std_logic_vector(9 downto 0);
    signal sumr_934 : std_logic_vector(9 downto 0);
    signal sumr_935 : std_logic_vector(9 downto 0);
    signal sumr_936 : std_logic_vector(9 downto 0);
    signal sumr_937 : std_logic_vector(9 downto 0);
    signal sumr_938 : std_logic_vector(9 downto 0);
    signal sumr_939 : std_logic_vector(9 downto 0);
    signal sumr_940 : std_logic_vector(9 downto 0);
    signal sumr_941 : std_logic_vector(9 downto 0);
    signal sumr_942 : std_logic_vector(9 downto 0);
    signal sumr_943 : std_logic_vector(9 downto 0);
    signal sumr_944 : std_logic_vector(9 downto 0);
    signal sumr_945 : std_logic_vector(9 downto 0);
    signal sumr_946 : std_logic_vector(9 downto 0);
    signal sumr_947 : std_logic_vector(9 downto 0);
    signal sumr_948 : std_logic_vector(9 downto 0);
    signal sumr_949 : std_logic_vector(9 downto 0);
    signal sumr_950 : std_logic_vector(9 downto 0);
    signal sumr_951 : std_logic_vector(9 downto 0);
    signal sumr_952 : std_logic_vector(9 downto 0);
    signal sumr_953 : std_logic_vector(9 downto 0);
    signal sumr_954 : std_logic_vector(9 downto 0);
    signal sumr_955 : std_logic_vector(9 downto 0);
    signal sumr_956 : std_logic_vector(9 downto 0);
    signal sumr_957 : std_logic_vector(9 downto 0);
    signal sumr_958 : std_logic_vector(9 downto 0);
    signal sumr_959 : std_logic_vector(9 downto 0);
    signal sumr_960 : std_logic_vector(9 downto 0);
    signal sumr_961 : std_logic_vector(9 downto 0);
    signal sumr_962 : std_logic_vector(9 downto 0);
    signal sumr_963 : std_logic_vector(9 downto 0);
    signal sumr_964 : std_logic_vector(9 downto 0);
    signal sumr_965 : std_logic_vector(9 downto 0);
    signal sumr_966 : std_logic_vector(9 downto 0);
    signal sumr_967 : std_logic_vector(9 downto 0);
    signal sumr_968 : std_logic_vector(9 downto 0);
    signal sumr_969 : std_logic_vector(9 downto 0);
    signal sumr_970 : std_logic_vector(9 downto 0);
    signal sumr_971 : std_logic_vector(9 downto 0);
    signal sumr_972 : std_logic_vector(9 downto 0);
    signal sumr_973 : std_logic_vector(9 downto 0);
    signal sumr_974 : std_logic_vector(9 downto 0);
    signal sumr_975 : std_logic_vector(9 downto 0);
    signal sumr_976 : std_logic_vector(9 downto 0);
    signal sumr_977 : std_logic_vector(9 downto 0);
    signal sumr_978 : std_logic_vector(9 downto 0);
    signal sumr_979 : std_logic_vector(9 downto 0);
    signal sumr_980 : std_logic_vector(9 downto 0);
    signal sumr_981 : std_logic_vector(9 downto 0);
    signal sumr_982 : std_logic_vector(9 downto 0);
    signal sumr_983 : std_logic_vector(9 downto 0);
    signal sumr_984 : std_logic_vector(9 downto 0);
    signal sumr_985 : std_logic_vector(9 downto 0);
    signal sumr_986 : std_logic_vector(9 downto 0);
    signal sumr_987 : std_logic_vector(9 downto 0);
    signal sumr_988 : std_logic_vector(9 downto 0);
    signal sumr_989 : std_logic_vector(9 downto 0);
    signal sumr_990 : std_logic_vector(9 downto 0);
    signal sumr_991 : std_logic_vector(9 downto 0);
    signal sumr_992 : std_logic_vector(9 downto 0);
    signal sumr_993 : std_logic_vector(9 downto 0);
    signal sumr_994 : std_logic_vector(9 downto 0);
    signal sumr_995 : std_logic_vector(9 downto 0);
    signal sumr_996 : std_logic_vector(9 downto 0);
    signal sumr_997 : std_logic_vector(9 downto 0);
    signal sumr_998 : std_logic_vector(9 downto 0);
    signal sumr_999 : std_logic_vector(9 downto 0);
    signal sumr_1000 : std_logic_vector(9 downto 0);
    signal sumr_1001 : std_logic_vector(9 downto 0);
    signal sumr_1002 : std_logic_vector(9 downto 0);
    signal sumr_1003 : std_logic_vector(9 downto 0);
    signal sumr_1004 : std_logic_vector(9 downto 0);
    signal sumr_1005 : std_logic_vector(9 downto 0);
    signal sumr_1006 : std_logic_vector(9 downto 0);
    signal sumr_1007 : std_logic_vector(9 downto 0);
    signal sumr_1008 : std_logic_vector(9 downto 0);
    signal sumr_1009 : std_logic_vector(9 downto 0);
    signal sumr_1010 : std_logic_vector(9 downto 0);
    signal sumr_1011 : std_logic_vector(9 downto 0);
    signal sumr_1012 : std_logic_vector(9 downto 0);
    signal sumr_1013 : std_logic_vector(9 downto 0);
    signal sumr_1014 : std_logic_vector(9 downto 0);
    signal sumr_1015 : std_logic_vector(9 downto 0);
    signal sumr_1016 : std_logic_vector(9 downto 0);
    signal sumr_1017 : std_logic_vector(9 downto 0);
    signal sumr_1018 : std_logic_vector(9 downto 0);
    signal sumr_1019 : std_logic_vector(9 downto 0);
    signal sumr_1020 : std_logic_vector(9 downto 0);
    signal sumr_1021 : std_logic_vector(9 downto 0);
    signal sumr_1022 : std_logic_vector(9 downto 0);
    signal sumr_1023 : std_logic_vector(9 downto 0);
begin

mulr_1_1<=a_1;
mulc_2_1 : entity work.gfmul
port map(
a=>a_2,
b=>"0000000010",
X=>mulr_2_1);

mulc_3_1 : entity work.gfmul
port map(
a=>a_3,
b=>"0000000100",
X=>mulr_3_1);

mulc_4_1 : entity work.gfmul
port map(
a=>a_4,
b=>"0000001000",
X=>mulr_4_1);

mulr_1_2<=a_1;
mulc_2_2 : entity work.gfmul
port map(
a=>a_2,
b=>"0000000100",
X=>mulr_2_2);

mulc_3_2 : entity work.gfmul
port map(
a=>a_3,
b=>"0000010000",
X=>mulr_3_2);

mulc_4_2 : entity work.gfmul
port map(
a=>a_4,
b=>"0001000000",
X=>mulr_4_2);

mulr_1_3<=a_1;
mulc_2_3 : entity work.gfmul
port map(
a=>a_2,
b=>"0000001000",
X=>mulr_2_3);

mulc_3_3 : entity work.gfmul
port map(
a=>a_3,
b=>"0001000000",
X=>mulr_3_3);

mulc_4_3 : entity work.gfmul
port map(
a=>a_4,
b=>"1000000000",
X=>mulr_4_3);

mulr_1_4<=a_1;
mulc_2_4 : entity work.gfmul
port map(
a=>a_2,
b=>"0000010000",
X=>mulr_2_4);

mulc_3_4 : entity work.gfmul
port map(
a=>a_3,
b=>"0100000000",
X=>mulr_3_4);

mulc_4_4 : entity work.gfmul
port map(
a=>a_4,
b=>"0000100100",
X=>mulr_4_4);

mulr_1_5<=a_1;
mulc_2_5 : entity work.gfmul
port map(
a=>a_2,
b=>"0000100000",
X=>mulr_2_5);

mulc_3_5 : entity work.gfmul
port map(
a=>a_3,
b=>"0000001001",
X=>mulr_3_5);

mulc_4_5 : entity work.gfmul
port map(
a=>a_4,
b=>"0100100000",
X=>mulr_4_5);

mulr_1_6<=a_1;
mulc_2_6 : entity work.gfmul
port map(
a=>a_2,
b=>"0001000000",
X=>mulr_2_6);

mulc_3_6 : entity work.gfmul
port map(
a=>a_3,
b=>"0000100100",
X=>mulr_3_6);

mulc_4_6 : entity work.gfmul
port map(
a=>a_4,
b=>"0100010010",
X=>mulr_4_6);

mulr_1_7<=a_1;
mulc_2_7 : entity work.gfmul
port map(
a=>a_2,
b=>"0010000000",
X=>mulr_2_7);

mulc_3_7 : entity work.gfmul
port map(
a=>a_3,
b=>"0010010000",
X=>mulr_3_7);

mulc_4_7 : entity work.gfmul
port map(
a=>a_4,
b=>"0010000010",
X=>mulr_4_7);

mulr_1_8<=a_1;
mulc_2_8 : entity work.gfmul
port map(
a=>a_2,
b=>"0100000000",
X=>mulr_2_8);

mulc_3_8 : entity work.gfmul
port map(
a=>a_3,
b=>"1001000000",
X=>mulr_3_8);

mulc_4_8 : entity work.gfmul
port map(
a=>a_4,
b=>"0000011001",
X=>mulr_4_8);

mulr_1_9<=a_1;
mulc_2_9 : entity work.gfmul
port map(
a=>a_2,
b=>"1000000000",
X=>mulr_2_9);

mulc_3_9 : entity work.gfmul
port map(
a=>a_3,
b=>"0100010010",
X=>mulr_3_9);

mulc_4_9 : entity work.gfmul
port map(
a=>a_4,
b=>"0011001000",
X=>mulr_4_9);

mulr_1_10<=a_1;
mulc_2_10 : entity work.gfmul
port map(
a=>a_2,
b=>"0000001001",
X=>mulr_2_10);

mulc_3_10 : entity work.gfmul
port map(
a=>a_3,
b=>"0001000001",
X=>mulr_3_10);

mulc_4_10 : entity work.gfmul
port map(
a=>a_4,
b=>"1001001001",
X=>mulr_4_10);

mulr_1_11<=a_1;
mulc_2_11 : entity work.gfmul
port map(
a=>a_2,
b=>"0000010010",
X=>mulr_2_11);

mulc_3_11 : entity work.gfmul
port map(
a=>a_3,
b=>"0100000100",
X=>mulr_3_11);

mulc_4_11 : entity work.gfmul
port map(
a=>a_4,
b=>"1001101100",
X=>mulr_4_11);

mulr_1_12<=a_1;
mulc_2_12 : entity work.gfmul
port map(
a=>a_2,
b=>"0000100100",
X=>mulr_2_12);

mulc_3_12 : entity work.gfmul
port map(
a=>a_3,
b=>"0000011001",
X=>mulr_3_12);

mulc_4_12 : entity work.gfmul
port map(
a=>a_4,
b=>"1101000100",
X=>mulr_4_12);

mulr_1_13<=a_1;
mulc_2_13 : entity work.gfmul
port map(
a=>a_2,
b=>"0001001000",
X=>mulr_2_13);

mulc_3_13 : entity work.gfmul
port map(
a=>a_3,
b=>"0001100100",
X=>mulr_3_13);

mulc_4_13 : entity work.gfmul
port map(
a=>a_4,
b=>"1000010110",
X=>mulr_4_13);

mulr_1_14<=a_1;
mulc_2_14 : entity work.gfmul
port map(
a=>a_2,
b=>"0010010000",
X=>mulr_2_14);

mulc_3_14 : entity work.gfmul
port map(
a=>a_3,
b=>"0110010000",
X=>mulr_3_14);

mulc_4_14 : entity work.gfmul
port map(
a=>a_4,
b=>"0010010100",
X=>mulr_4_14);

mulr_1_15<=a_1;
mulc_2_15 : entity work.gfmul
port map(
a=>a_2,
b=>"0100100000",
X=>mulr_2_15);

mulc_3_15 : entity work.gfmul
port map(
a=>a_3,
b=>"1001001001",
X=>mulr_3_15);

mulc_4_15 : entity work.gfmul
port map(
a=>a_4,
b=>"0010101001",
X=>mulr_4_15);

mulr_1_16<=a_1;
mulc_2_16 : entity work.gfmul
port map(
a=>a_2,
b=>"1001000000",
X=>mulr_2_16);

mulc_3_16 : entity work.gfmul
port map(
a=>a_3,
b=>"0100110110",
X=>mulr_3_16);

mulc_4_16 : entity work.gfmul
port map(
a=>a_4,
b=>"0101000001",
X=>mulr_4_16);

mulr_1_17<=a_1;
mulc_2_17 : entity work.gfmul
port map(
a=>a_2,
b=>"0010001001",
X=>mulr_2_17);

mulc_3_17 : entity work.gfmul
port map(
a=>a_3,
b=>"0011010001",
X=>mulr_3_17);

mulc_4_17 : entity work.gfmul
port map(
a=>a_4,
b=>"1000011010",
X=>mulr_4_17);

mulr_1_18<=a_1;
mulc_2_18 : entity work.gfmul
port map(
a=>a_2,
b=>"0100010010",
X=>mulr_2_18);

mulc_3_18 : entity work.gfmul
port map(
a=>a_3,
b=>"1101000100",
X=>mulr_3_18);

mulc_4_18 : entity work.gfmul
port map(
a=>a_4,
b=>"0011110100",
X=>mulr_4_18);

mulr_1_19<=a_1;
mulc_2_19 : entity work.gfmul
port map(
a=>a_2,
b=>"1000100100",
X=>mulr_2_19);

mulc_3_19 : entity work.gfmul
port map(
a=>a_3,
b=>"0100001011",
X=>mulr_3_19);

mulc_4_19 : entity work.gfmul
port map(
a=>a_4,
b=>"1110101001",
X=>mulr_4_19);

mulr_1_20<=a_1;
mulc_2_20 : entity work.gfmul
port map(
a=>a_2,
b=>"0001000001",
X=>mulr_2_20);

mulc_3_20 : entity work.gfmul
port map(
a=>a_3,
b=>"0000100101",
X=>mulr_3_20);

mulc_4_20 : entity work.gfmul
port map(
a=>a_4,
b=>"0101110111",
X=>mulr_4_20);

mulr_1_21<=a_1;
mulc_2_21 : entity work.gfmul
port map(
a=>a_2,
b=>"0010000010",
X=>mulr_2_21);

mulc_3_21 : entity work.gfmul
port map(
a=>a_3,
b=>"0010010100",
X=>mulr_3_21);

mulc_4_21 : entity work.gfmul
port map(
a=>a_4,
b=>"1110101010",
X=>mulr_4_21);

mulr_1_22<=a_1;
mulc_2_22 : entity work.gfmul
port map(
a=>a_2,
b=>"0100000100",
X=>mulr_2_22);

mulc_3_22 : entity work.gfmul
port map(
a=>a_3,
b=>"1001010000",
X=>mulr_3_22);

mulc_4_22 : entity work.gfmul
port map(
a=>a_4,
b=>"0101101111",
X=>mulr_4_22);

mulr_1_23<=a_1;
mulc_2_23 : entity work.gfmul
port map(
a=>a_2,
b=>"1000001000",
X=>mulr_2_23);

mulc_3_23 : entity work.gfmul
port map(
a=>a_3,
b=>"0101010010",
X=>mulr_3_23);

mulc_4_23 : entity work.gfmul
port map(
a=>a_4,
b=>"1101101010",
X=>mulr_4_23);

mulr_1_24<=a_1;
mulc_2_24 : entity work.gfmul
port map(
a=>a_2,
b=>"0000011001",
X=>mulr_2_24);

mulc_3_24 : entity work.gfmul
port map(
a=>a_3,
b=>"0101000001",
X=>mulr_3_24);

mulc_4_24 : entity work.gfmul
port map(
a=>a_4,
b=>"1101100110",
X=>mulr_4_24);

mulr_1_25<=a_1;
mulc_2_25 : entity work.gfmul
port map(
a=>a_2,
b=>"0000110010",
X=>mulr_2_25);

mulc_3_25 : entity work.gfmul
port map(
a=>a_3,
b=>"0100001101",
X=>mulr_3_25);

mulc_4_25 : entity work.gfmul
port map(
a=>a_4,
b=>"1100000110",
X=>mulr_4_25);

mulr_1_26<=a_1;
mulc_2_26 : entity work.gfmul
port map(
a=>a_2,
b=>"0001100100",
X=>mulr_2_26);

mulc_3_26 : entity work.gfmul
port map(
a=>a_3,
b=>"0000111101",
X=>mulr_3_26);

mulc_4_26 : entity work.gfmul
port map(
a=>a_4,
b=>"0000000110",
X=>mulr_4_26);

mulr_1_27<=a_1;
mulc_2_27 : entity work.gfmul
port map(
a=>a_2,
b=>"0011001000",
X=>mulr_2_27);

mulc_3_27 : entity work.gfmul
port map(
a=>a_3,
b=>"0011110100",
X=>mulr_3_27);

mulc_4_27 : entity work.gfmul
port map(
a=>a_4,
b=>"0000110000",
X=>mulr_4_27);

mulr_1_28<=a_1;
mulc_2_28 : entity work.gfmul
port map(
a=>a_2,
b=>"0110010000",
X=>mulr_2_28);

mulc_3_28 : entity work.gfmul
port map(
a=>a_3,
b=>"1111010000",
X=>mulr_3_28);

mulc_4_28 : entity work.gfmul
port map(
a=>a_4,
b=>"0110000000",
X=>mulr_4_28);

mulr_1_29<=a_1;
mulc_2_29 : entity work.gfmul
port map(
a=>a_2,
b=>"1100100000",
X=>mulr_2_29);

mulc_3_29 : entity work.gfmul
port map(
a=>a_3,
b=>"1101011011",
X=>mulr_3_29);

mulc_4_29 : entity work.gfmul
port map(
a=>a_4,
b=>"0000011011",
X=>mulr_4_29);

mulr_1_30<=a_1;
mulc_2_30 : entity work.gfmul
port map(
a=>a_2,
b=>"1001001001",
X=>mulr_2_30);

mulc_3_30 : entity work.gfmul
port map(
a=>a_3,
b=>"0101110111",
X=>mulr_3_30);

mulc_4_30 : entity work.gfmul
port map(
a=>a_4,
b=>"0011011000",
X=>mulr_4_30);

mulr_1_31<=a_1;
mulc_2_31 : entity work.gfmul
port map(
a=>a_2,
b=>"0010011011",
X=>mulr_2_31);

mulc_3_31 : entity work.gfmul
port map(
a=>a_3,
b=>"0111010101",
X=>mulr_3_31);

mulc_4_31 : entity work.gfmul
port map(
a=>a_4,
b=>"1011001001",
X=>mulr_4_31);

mulr_1_32<=a_1;
mulc_2_32 : entity work.gfmul
port map(
a=>a_2,
b=>"0100110110",
X=>mulr_2_32);

mulc_3_32 : entity work.gfmul
port map(
a=>a_3,
b=>"1101011101",
X=>mulr_3_32);

mulc_4_32 : entity work.gfmul
port map(
a=>a_4,
b=>"1001100101",
X=>mulr_4_32);

mulr_1_33<=a_1;
mulc_2_33 : entity work.gfmul
port map(
a=>a_2,
b=>"1001101100",
X=>mulr_2_33);

mulc_3_33 : entity work.gfmul
port map(
a=>a_3,
b=>"0101101111",
X=>mulr_3_33);

mulc_4_33 : entity work.gfmul
port map(
a=>a_4,
b=>"1100001100",
X=>mulr_4_33);

mulr_1_34<=a_1;
mulc_2_34 : entity work.gfmul
port map(
a=>a_2,
b=>"0011010001",
X=>mulr_2_34);

mulc_3_34 : entity work.gfmul
port map(
a=>a_3,
b=>"0110110101",
X=>mulr_3_34);

mulc_4_34 : entity work.gfmul
port map(
a=>a_4,
b=>"0001010110",
X=>mulr_4_34);

mulr_1_35<=a_1;
mulc_2_35 : entity work.gfmul
port map(
a=>a_2,
b=>"0110100010",
X=>mulr_2_35);

mulc_3_35 : entity work.gfmul
port map(
a=>a_3,
b=>"1011011101",
X=>mulr_3_35);

mulc_4_35 : entity work.gfmul
port map(
a=>a_4,
b=>"1010110000",
X=>mulr_4_35);

mulr_1_36<=a_1;
mulc_2_36 : entity work.gfmul
port map(
a=>a_2,
b=>"1101000100",
X=>mulr_2_36);

mulc_3_36 : entity work.gfmul
port map(
a=>a_3,
b=>"1101100110",
X=>mulr_3_36);

mulc_4_36 : entity work.gfmul
port map(
a=>a_4,
b=>"0110101101",
X=>mulr_4_36);

mulr_1_37<=a_1;
mulc_2_37 : entity work.gfmul
port map(
a=>a_2,
b=>"1010000001",
X=>mulr_2_37);

mulc_3_37 : entity work.gfmul
port map(
a=>a_3,
b=>"0110000011",
X=>mulr_3_37);

mulc_4_37 : entity work.gfmul
port map(
a=>a_4,
b=>"0101110011",
X=>mulr_4_37);

mulr_1_38<=a_1;
mulc_2_38 : entity work.gfmul
port map(
a=>a_2,
b=>"0100001011",
X=>mulr_2_38);

mulc_3_38 : entity work.gfmul
port map(
a=>a_3,
b=>"1000000101",
X=>mulr_3_38);

mulc_4_38 : entity work.gfmul
port map(
a=>a_4,
b=>"1110001010",
X=>mulr_4_38);

mulr_1_39<=a_1;
mulc_2_39 : entity work.gfmul
port map(
a=>a_2,
b=>"1000010110",
X=>mulr_2_39);

mulc_3_39 : entity work.gfmul
port map(
a=>a_3,
b=>"0000000110",
X=>mulr_3_39);

mulc_4_39 : entity work.gfmul
port map(
a=>a_4,
b=>"0001101111",
X=>mulr_4_39);

mulr_1_40<=a_1;
mulc_2_40 : entity work.gfmul
port map(
a=>a_2,
b=>"0000100101",
X=>mulr_2_40);

mulc_3_40 : entity work.gfmul
port map(
a=>a_3,
b=>"0000011000",
X=>mulr_3_40);

mulc_4_40 : entity work.gfmul
port map(
a=>a_4,
b=>"1101111000",
X=>mulr_4_40);

mulr_1_41<=a_1;
mulc_2_41 : entity work.gfmul
port map(
a=>a_2,
b=>"0001001010",
X=>mulr_2_41);

mulc_3_41 : entity work.gfmul
port map(
a=>a_3,
b=>"0001100000",
X=>mulr_3_41);

mulc_4_41 : entity work.gfmul
port map(
a=>a_4,
b=>"1111110110",
X=>mulr_4_41);

mulr_1_42<=a_1;
mulc_2_42 : entity work.gfmul
port map(
a=>a_2,
b=>"0010010100",
X=>mulr_2_42);

mulc_3_42 : entity work.gfmul
port map(
a=>a_3,
b=>"0110000000",
X=>mulr_3_42);

mulc_4_42 : entity work.gfmul
port map(
a=>a_4,
b=>"1110001111",
X=>mulr_4_42);

mulr_1_43<=a_1;
mulc_2_43 : entity work.gfmul
port map(
a=>a_2,
b=>"0100101000",
X=>mulr_2_43);

mulc_3_43 : entity work.gfmul
port map(
a=>a_3,
b=>"1000001001",
X=>mulr_3_43);

mulc_4_43 : entity work.gfmul
port map(
a=>a_4,
b=>"0001000111",
X=>mulr_4_43);

mulr_1_44<=a_1;
mulc_2_44 : entity work.gfmul
port map(
a=>a_2,
b=>"1001010000",
X=>mulr_2_44);

mulc_3_44 : entity work.gfmul
port map(
a=>a_3,
b=>"0000110110",
X=>mulr_3_44);

mulc_4_44 : entity work.gfmul
port map(
a=>a_4,
b=>"1000111000",
X=>mulr_4_44);

mulr_1_45<=a_1;
mulc_2_45 : entity work.gfmul
port map(
a=>a_2,
b=>"0010101001",
X=>mulr_2_45);

mulc_3_45 : entity work.gfmul
port map(
a=>a_3,
b=>"0011011000",
X=>mulr_3_45);

mulc_4_45 : entity work.gfmul
port map(
a=>a_4,
b=>"0111100100",
X=>mulr_4_45);

mulr_1_46<=a_1;
mulc_2_46 : entity work.gfmul
port map(
a=>a_2,
b=>"0101010010",
X=>mulr_2_46);

mulc_3_46 : entity work.gfmul
port map(
a=>a_3,
b=>"1101100000",
X=>mulr_3_46);

mulc_4_46 : entity work.gfmul
port map(
a=>a_4,
b=>"1100111011",
X=>mulr_4_46);

mulr_1_47<=a_1;
mulc_2_47 : entity work.gfmul
port map(
a=>a_2,
b=>"1010100100",
X=>mulr_2_47);

mulc_3_47 : entity work.gfmul
port map(
a=>a_3,
b=>"0110011011",
X=>mulr_3_47);

mulc_4_47 : entity work.gfmul
port map(
a=>a_4,
b=>"0111101110",
X=>mulr_4_47);

mulr_1_48<=a_1;
mulc_2_48 : entity work.gfmul
port map(
a=>a_2,
b=>"0101000001",
X=>mulr_2_48);

mulc_3_48 : entity work.gfmul
port map(
a=>a_3,
b=>"1001100101",
X=>mulr_3_48);

mulc_4_48 : entity work.gfmul
port map(
a=>a_4,
b=>"1101101011",
X=>mulr_4_48);

mulr_1_49<=a_1;
mulc_2_49 : entity work.gfmul
port map(
a=>a_2,
b=>"1010000010",
X=>mulr_2_49);

mulc_3_49 : entity work.gfmul
port map(
a=>a_3,
b=>"0110000110",
X=>mulr_3_49);

mulc_4_49 : entity work.gfmul
port map(
a=>a_4,
b=>"1101101110",
X=>mulr_4_49);

mulr_1_50<=a_1;
mulc_2_50 : entity work.gfmul
port map(
a=>a_2,
b=>"0100001101",
X=>mulr_2_50);

mulc_3_50 : entity work.gfmul
port map(
a=>a_3,
b=>"1000010001",
X=>mulr_3_50);

mulc_4_50 : entity work.gfmul
port map(
a=>a_4,
b=>"1101000110",
X=>mulr_4_50);

mulr_1_51<=a_1;
mulc_2_51 : entity work.gfmul
port map(
a=>a_2,
b=>"1000011010",
X=>mulr_2_51);

mulc_3_51 : entity work.gfmul
port map(
a=>a_3,
b=>"0001010110",
X=>mulr_3_51);

mulc_4_51 : entity work.gfmul
port map(
a=>a_4,
b=>"1000000110",
X=>mulr_4_51);

mulr_1_52<=a_1;
mulc_2_52 : entity work.gfmul
port map(
a=>a_2,
b=>"0000111101",
X=>mulr_2_52);

mulc_3_52 : entity work.gfmul
port map(
a=>a_3,
b=>"0101011000",
X=>mulr_3_52);

mulc_4_52 : entity work.gfmul
port map(
a=>a_4,
b=>"0000010100",
X=>mulr_4_52);

mulr_1_53<=a_1;
mulc_2_53 : entity work.gfmul
port map(
a=>a_2,
b=>"0001111010",
X=>mulr_2_53);

mulc_3_53 : entity work.gfmul
port map(
a=>a_3,
b=>"0101101001",
X=>mulr_3_53);

mulc_4_53 : entity work.gfmul
port map(
a=>a_4,
b=>"0010100000",
X=>mulr_4_53);

mulr_1_54<=a_1;
mulc_2_54 : entity work.gfmul
port map(
a=>a_2,
b=>"0011110100",
X=>mulr_2_54);

mulc_3_54 : entity work.gfmul
port map(
a=>a_3,
b=>"0110101101",
X=>mulr_3_54);

mulc_4_54 : entity work.gfmul
port map(
a=>a_4,
b=>"0100001001",
X=>mulr_4_54);

mulr_1_55<=a_1;
mulc_2_55 : entity work.gfmul
port map(
a=>a_2,
b=>"0111101000",
X=>mulr_2_55);

mulc_3_55 : entity work.gfmul
port map(
a=>a_3,
b=>"1010111101",
X=>mulr_3_55);

mulc_4_55 : entity work.gfmul
port map(
a=>a_4,
b=>"0001011010",
X=>mulr_4_55);

mulr_1_56<=a_1;
mulc_2_56 : entity work.gfmul
port map(
a=>a_2,
b=>"1111010000",
X=>mulr_2_56);

mulc_3_56 : entity work.gfmul
port map(
a=>a_3,
b=>"1011100110",
X=>mulr_3_56);

mulc_4_56 : entity work.gfmul
port map(
a=>a_4,
b=>"1011010000",
X=>mulr_4_56);

mulr_1_57<=a_1;
mulc_2_57 : entity work.gfmul
port map(
a=>a_2,
b=>"1110101001",
X=>mulr_2_57);

mulc_3_57 : entity work.gfmul
port map(
a=>a_3,
b=>"1110001010",
X=>mulr_3_57);

mulc_4_57 : entity work.gfmul
port map(
a=>a_4,
b=>"1010101101",
X=>mulr_4_57);

mulr_1_58<=a_1;
mulc_2_58 : entity work.gfmul
port map(
a=>a_2,
b=>"1101011011",
X=>mulr_2_58);

mulc_3_58 : entity work.gfmul
port map(
a=>a_3,
b=>"1000110011",
X=>mulr_3_58);

mulc_4_58 : entity work.gfmul
port map(
a=>a_4,
b=>"0101000101",
X=>mulr_4_58);

mulr_1_59<=a_1;
mulc_2_59 : entity work.gfmul
port map(
a=>a_2,
b=>"1010111111",
X=>mulr_2_59);

mulc_3_59 : entity work.gfmul
port map(
a=>a_3,
b=>"0011011110",
X=>mulr_3_59);

mulc_4_59 : entity work.gfmul
port map(
a=>a_4,
b=>"1000111010",
X=>mulr_4_59);

mulr_1_60<=a_1;
mulc_2_60 : entity work.gfmul
port map(
a=>a_2,
b=>"0101110111",
X=>mulr_2_60);

mulc_3_60 : entity work.gfmul
port map(
a=>a_3,
b=>"1101111000",
X=>mulr_3_60);

mulc_4_60 : entity work.gfmul
port map(
a=>a_4,
b=>"0111110100",
X=>mulr_4_60);

mulr_1_61<=a_1;
mulc_2_61 : entity work.gfmul
port map(
a=>a_2,
b=>"1011101110",
X=>mulr_2_61);

mulc_3_61 : entity work.gfmul
port map(
a=>a_3,
b=>"0111111011",
X=>mulr_3_61);

mulc_4_61 : entity work.gfmul
port map(
a=>a_4,
b=>"1110111011",
X=>mulr_4_61);

mulr_1_62<=a_1;
mulc_2_62 : entity work.gfmul
port map(
a=>a_2,
b=>"0111010101",
X=>mulr_2_62);

mulc_3_62 : entity work.gfmul
port map(
a=>a_3,
b=>"1111100101",
X=>mulr_3_62);

mulc_4_62 : entity work.gfmul
port map(
a=>a_4,
b=>"0111100111",
X=>mulr_4_62);

mulr_1_63<=a_1;
mulc_2_63 : entity work.gfmul
port map(
a=>a_2,
b=>"1110101010",
X=>mulr_2_63);

mulc_3_63 : entity work.gfmul
port map(
a=>a_3,
b=>"1110001111",
X=>mulr_3_63);

mulc_4_63 : entity work.gfmul
port map(
a=>a_4,
b=>"1100100011",
X=>mulr_4_63);

mulr_1_64<=a_1;
mulc_2_64 : entity work.gfmul
port map(
a=>a_2,
b=>"1101011101",
X=>mulr_2_64);

mulc_3_64 : entity work.gfmul
port map(
a=>a_3,
b=>"1000100111",
X=>mulr_3_64);

mulc_4_64 : entity work.gfmul
port map(
a=>a_4,
b=>"0100101110",
X=>mulr_4_64);

mulr_1_65<=a_1;
mulc_2_65 : entity work.gfmul
port map(
a=>a_2,
b=>"1010110011",
X=>mulr_2_65);

mulc_3_65 : entity work.gfmul
port map(
a=>a_3,
b=>"0010001110",
X=>mulr_3_65);

mulc_4_65 : entity work.gfmul
port map(
a=>a_4,
b=>"0101100010",
X=>mulr_4_65);

mulr_1_66<=a_1;
mulc_2_66 : entity work.gfmul
port map(
a=>a_2,
b=>"0101101111",
X=>mulr_2_66);

mulc_3_66 : entity work.gfmul
port map(
a=>a_3,
b=>"1000111000",
X=>mulr_3_66);

mulc_4_66 : entity work.gfmul
port map(
a=>a_4,
b=>"1100000010",
X=>mulr_4_66);

mulr_1_67<=a_1;
mulc_2_67 : entity work.gfmul
port map(
a=>a_2,
b=>"1011011110",
X=>mulr_2_67);

mulc_3_67 : entity work.gfmul
port map(
a=>a_3,
b=>"0011110010",
X=>mulr_3_67);

mulc_4_67 : entity work.gfmul
port map(
a=>a_4,
b=>"0000100110",
X=>mulr_4_67);

mulr_1_68<=a_1;
mulc_2_68 : entity work.gfmul
port map(
a=>a_2,
b=>"0110110101",
X=>mulr_2_68);

mulc_3_68 : entity work.gfmul
port map(
a=>a_3,
b=>"1111001000",
X=>mulr_3_68);

mulc_4_68 : entity work.gfmul
port map(
a=>a_4,
b=>"0100110000",
X=>mulr_4_68);

mulr_1_69<=a_1;
mulc_2_69 : entity work.gfmul
port map(
a=>a_2,
b=>"1101101010",
X=>mulr_2_69);

mulc_3_69 : entity work.gfmul
port map(
a=>a_3,
b=>"1100111011",
X=>mulr_3_69);

mulc_4_69 : entity work.gfmul
port map(
a=>a_4,
b=>"0110010010",
X=>mulr_4_69);

mulr_1_70<=a_1;
mulc_2_70 : entity work.gfmul
port map(
a=>a_2,
b=>"1011011101",
X=>mulr_2_70);

mulc_3_70 : entity work.gfmul
port map(
a=>a_3,
b=>"0011110111",
X=>mulr_3_70);

mulc_4_70 : entity work.gfmul
port map(
a=>a_4,
b=>"0010001011",
X=>mulr_4_70);

mulr_1_71<=a_1;
mulc_2_71 : entity work.gfmul
port map(
a=>a_2,
b=>"0110110011",
X=>mulr_2_71);

mulc_3_71 : entity work.gfmul
port map(
a=>a_3,
b=>"1111011100",
X=>mulr_3_71);

mulc_4_71 : entity work.gfmul
port map(
a=>a_4,
b=>"0001010001",
X=>mulr_4_71);

mulr_1_72<=a_1;
mulc_2_72 : entity work.gfmul
port map(
a=>a_2,
b=>"1101100110",
X=>mulr_2_72);

mulc_3_72 : entity work.gfmul
port map(
a=>a_3,
b=>"1101101011",
X=>mulr_3_72);

mulc_4_72 : entity work.gfmul
port map(
a=>a_4,
b=>"1010001000",
X=>mulr_4_72);

mulr_1_73<=a_1;
mulc_2_73 : entity work.gfmul
port map(
a=>a_2,
b=>"1011000101",
X=>mulr_2_73);

mulc_3_73 : entity work.gfmul
port map(
a=>a_3,
b=>"0110110111",
X=>mulr_3_73);

mulc_4_73 : entity work.gfmul
port map(
a=>a_4,
b=>"0001101101",
X=>mulr_4_73);

mulr_1_74<=a_1;
mulc_2_74 : entity work.gfmul
port map(
a=>a_2,
b=>"0110000011",
X=>mulr_2_74);

mulc_3_74 : entity work.gfmul
port map(
a=>a_3,
b=>"1011010101",
X=>mulr_3_74);

mulc_4_74 : entity work.gfmul
port map(
a=>a_4,
b=>"1101101000",
X=>mulr_4_74);

mulr_1_75<=a_1;
mulc_2_75 : entity work.gfmul
port map(
a=>a_2,
b=>"1100000110",
X=>mulr_2_75);

mulc_3_75 : entity work.gfmul
port map(
a=>a_3,
b=>"1101000110",
X=>mulr_3_75);

mulc_4_75 : entity work.gfmul
port map(
a=>a_4,
b=>"1101110110",
X=>mulr_4_75);

mulr_1_76<=a_1;
mulc_2_76 : entity work.gfmul
port map(
a=>a_2,
b=>"1000000101",
X=>mulr_2_76);

mulc_3_76 : entity work.gfmul
port map(
a=>a_3,
b=>"0100000011",
X=>mulr_3_76);

mulc_4_76 : entity work.gfmul
port map(
a=>a_4,
b=>"1110000110",
X=>mulr_4_76);

mulr_1_77<=a_1;
mulc_2_77 : entity work.gfmul
port map(
a=>a_2,
b=>"0000000011",
X=>mulr_2_77);

mulc_3_77 : entity work.gfmul
port map(
a=>a_3,
b=>"0000000101",
X=>mulr_3_77);

mulc_4_77 : entity work.gfmul
port map(
a=>a_4,
b=>"0000001111",
X=>mulr_4_77);

mulr_1_78<=a_1;
mulc_2_78 : entity work.gfmul
port map(
a=>a_2,
b=>"0000000110",
X=>mulr_2_78);

mulc_3_78 : entity work.gfmul
port map(
a=>a_3,
b=>"0000010100",
X=>mulr_3_78);

mulc_4_78 : entity work.gfmul
port map(
a=>a_4,
b=>"0001111000",
X=>mulr_4_78);

mulr_1_79<=a_1;
mulc_2_79 : entity work.gfmul
port map(
a=>a_2,
b=>"0000001100",
X=>mulr_2_79);

mulc_3_79 : entity work.gfmul
port map(
a=>a_3,
b=>"0001010000",
X=>mulr_3_79);

mulc_4_79 : entity work.gfmul
port map(
a=>a_4,
b=>"1111000000",
X=>mulr_4_79);

mulr_1_80<=a_1;
mulc_2_80 : entity work.gfmul
port map(
a=>a_2,
b=>"0000011000",
X=>mulr_2_80);

mulc_3_80 : entity work.gfmul
port map(
a=>a_3,
b=>"0101000000",
X=>mulr_3_80);

mulc_4_80 : entity work.gfmul
port map(
a=>a_4,
b=>"1000111111",
X=>mulr_4_80);

mulr_1_81<=a_1;
mulc_2_81 : entity work.gfmul
port map(
a=>a_2,
b=>"0000110000",
X=>mulr_2_81);

mulc_3_81 : entity work.gfmul
port map(
a=>a_3,
b=>"0100001001",
X=>mulr_3_81);

mulc_4_81 : entity work.gfmul
port map(
a=>a_4,
b=>"0111011100",
X=>mulr_4_81);

mulr_1_82<=a_1;
mulc_2_82 : entity work.gfmul
port map(
a=>a_2,
b=>"0001100000",
X=>mulr_2_82);

mulc_3_82 : entity work.gfmul
port map(
a=>a_3,
b=>"0000101101",
X=>mulr_3_82);

mulc_4_82 : entity work.gfmul
port map(
a=>a_4,
b=>"1011111011",
X=>mulr_4_82);

mulr_1_83<=a_1;
mulc_2_83 : entity work.gfmul
port map(
a=>a_2,
b=>"0011000000",
X=>mulr_2_83);

mulc_3_83 : entity work.gfmul
port map(
a=>a_3,
b=>"0010110100",
X=>mulr_3_83);

mulc_4_83 : entity work.gfmul
port map(
a=>a_4,
b=>"1111110101",
X=>mulr_4_83);

mulr_1_84<=a_1;
mulc_2_84 : entity work.gfmul
port map(
a=>a_2,
b=>"0110000000",
X=>mulr_2_84);

mulc_3_84 : entity work.gfmul
port map(
a=>a_3,
b=>"1011010000",
X=>mulr_3_84);

mulc_4_84 : entity work.gfmul
port map(
a=>a_4,
b=>"1110010111",
X=>mulr_4_84);

mulr_1_85<=a_1;
mulc_2_85 : entity work.gfmul
port map(
a=>a_2,
b=>"1100000000",
X=>mulr_2_85);

mulc_3_85 : entity work.gfmul
port map(
a=>a_3,
b=>"1101010010",
X=>mulr_3_85);

mulc_4_85 : entity work.gfmul
port map(
a=>a_4,
b=>"0010000111",
X=>mulr_4_85);

mulr_1_86<=a_1;
mulc_2_86 : entity work.gfmul
port map(
a=>a_2,
b=>"1000001001",
X=>mulr_2_86);

mulc_3_86 : entity work.gfmul
port map(
a=>a_3,
b=>"0101010011",
X=>mulr_3_86);

mulc_4_86 : entity work.gfmul
port map(
a=>a_4,
b=>"0000110001",
X=>mulr_4_86);

mulr_1_87<=a_1;
mulc_2_87 : entity work.gfmul
port map(
a=>a_2,
b=>"0000011011",
X=>mulr_2_87);

mulc_3_87 : entity work.gfmul
port map(
a=>a_3,
b=>"0101000101",
X=>mulr_3_87);

mulc_4_87 : entity work.gfmul
port map(
a=>a_4,
b=>"0110001000",
X=>mulr_4_87);

mulr_1_88<=a_1;
mulc_2_88 : entity work.gfmul
port map(
a=>a_2,
b=>"0000110110",
X=>mulr_2_88);

mulc_3_88 : entity work.gfmul
port map(
a=>a_3,
b=>"0100011101",
X=>mulr_3_88);

mulc_4_88 : entity work.gfmul
port map(
a=>a_4,
b=>"0001011011",
X=>mulr_4_88);

mulr_1_89<=a_1;
mulc_2_89 : entity work.gfmul
port map(
a=>a_2,
b=>"0001101100",
X=>mulr_2_89);

mulc_3_89 : entity work.gfmul
port map(
a=>a_3,
b=>"0001111101",
X=>mulr_3_89);

mulc_4_89 : entity work.gfmul
port map(
a=>a_4,
b=>"1011011000",
X=>mulr_4_89);

mulr_1_90<=a_1;
mulc_2_90 : entity work.gfmul
port map(
a=>a_2,
b=>"0011011000",
X=>mulr_2_90);

mulc_3_90 : entity work.gfmul
port map(
a=>a_3,
b=>"0111110100",
X=>mulr_3_90);

mulc_4_90 : entity work.gfmul
port map(
a=>a_4,
b=>"1011101101",
X=>mulr_4_90);

mulr_1_91<=a_1;
mulc_2_91 : entity work.gfmul
port map(
a=>a_2,
b=>"0110110000",
X=>mulr_2_91);

mulc_3_91 : entity work.gfmul
port map(
a=>a_3,
b=>"1111011001",
X=>mulr_3_91);

mulc_4_91 : entity work.gfmul
port map(
a=>a_4,
b=>"1101000101",
X=>mulr_4_91);

mulr_1_92<=a_1;
mulc_2_92 : entity work.gfmul
port map(
a=>a_2,
b=>"1101100000",
X=>mulr_2_92);

mulc_3_92 : entity work.gfmul
port map(
a=>a_3,
b=>"1101111111",
X=>mulr_3_92);

mulc_4_92 : entity work.gfmul
port map(
a=>a_4,
b=>"1000011110",
X=>mulr_4_92);

mulr_1_93<=a_1;
mulc_2_93 : entity work.gfmul
port map(
a=>a_2,
b=>"1011001001",
X=>mulr_2_93);

mulc_3_93 : entity work.gfmul
port map(
a=>a_3,
b=>"0111100111",
X=>mulr_3_93);

mulc_4_93 : entity work.gfmul
port map(
a=>a_4,
b=>"0011010100",
X=>mulr_4_93);

mulr_1_94<=a_1;
mulc_2_94 : entity work.gfmul
port map(
a=>a_2,
b=>"0110011011",
X=>mulr_2_94);

mulc_3_94 : entity work.gfmul
port map(
a=>a_3,
b=>"1110010101",
X=>mulr_3_94);

mulc_4_94 : entity work.gfmul
port map(
a=>a_4,
b=>"1010101001",
X=>mulr_4_94);

mulr_1_95<=a_1;
mulc_2_95 : entity work.gfmul
port map(
a=>a_2,
b=>"1100110110",
X=>mulr_2_95);

mulc_3_95 : entity work.gfmul
port map(
a=>a_3,
b=>"1001001111",
X=>mulr_3_95);

mulc_4_95 : entity work.gfmul
port map(
a=>a_4,
b=>"0101100101",
X=>mulr_4_95);

mulr_1_96<=a_1;
mulc_2_96 : entity work.gfmul
port map(
a=>a_2,
b=>"1001100101",
X=>mulr_2_96);

mulc_3_96 : entity work.gfmul
port map(
a=>a_3,
b=>"0100101110",
X=>mulr_3_96);

mulc_4_96 : entity work.gfmul
port map(
a=>a_4,
b=>"1100111010",
X=>mulr_4_96);

mulr_1_97<=a_1;
mulc_2_97 : entity work.gfmul
port map(
a=>a_2,
b=>"0011000011",
X=>mulr_2_97);

mulc_3_97 : entity work.gfmul
port map(
a=>a_3,
b=>"0010110001",
X=>mulr_3_97);

mulc_4_97 : entity work.gfmul
port map(
a=>a_4,
b=>"0111100110",
X=>mulr_4_97);

mulr_1_98<=a_1;
mulc_2_98 : entity work.gfmul
port map(
a=>a_2,
b=>"0110000110",
X=>mulr_2_98);

mulc_3_98 : entity work.gfmul
port map(
a=>a_3,
b=>"1011000100",
X=>mulr_3_98);

mulc_4_98 : entity work.gfmul
port map(
a=>a_4,
b=>"1100101011",
X=>mulr_4_98);

mulr_1_99<=a_1;
mulc_2_99 : entity work.gfmul
port map(
a=>a_2,
b=>"1100001100",
X=>mulr_2_99);

mulc_3_99 : entity work.gfmul
port map(
a=>a_3,
b=>"1100000010",
X=>mulr_3_99);

mulc_4_99 : entity work.gfmul
port map(
a=>a_4,
b=>"0101101110",
X=>mulr_4_99);

mulr_1_100<=a_1;
mulc_2_100 : entity work.gfmul
port map(
a=>a_2,
b=>"1000010001",
X=>mulr_2_100);

mulc_3_100 : entity work.gfmul
port map(
a=>a_3,
b=>"0000010011",
X=>mulr_3_100);

mulc_4_100 : entity work.gfmul
port map(
a=>a_4,
b=>"1101100010",
X=>mulr_4_100);

mulr_1_101<=a_1;
mulc_2_101 : entity work.gfmul
port map(
a=>a_2,
b=>"0000101011",
X=>mulr_2_101);

mulc_3_101 : entity work.gfmul
port map(
a=>a_3,
b=>"0001001100",
X=>mulr_3_101);

mulc_4_101 : entity work.gfmul
port map(
a=>a_4,
b=>"1100100110",
X=>mulr_4_101);

mulr_1_102<=a_1;
mulc_2_102 : entity work.gfmul
port map(
a=>a_2,
b=>"0001010110",
X=>mulr_2_102);

mulc_3_102 : entity work.gfmul
port map(
a=>a_3,
b=>"0100110000",
X=>mulr_3_102);

mulc_4_102 : entity work.gfmul
port map(
a=>a_4,
b=>"0100000110",
X=>mulr_4_102);

mulr_1_103<=a_1;
mulc_2_103 : entity work.gfmul
port map(
a=>a_2,
b=>"0010101100",
X=>mulr_2_103);

mulc_3_103 : entity work.gfmul
port map(
a=>a_3,
b=>"0011001001",
X=>mulr_3_103);

mulc_4_103 : entity work.gfmul
port map(
a=>a_4,
b=>"0000100010",
X=>mulr_4_103);

mulr_1_104<=a_1;
mulc_2_104 : entity work.gfmul
port map(
a=>a_2,
b=>"0101011000",
X=>mulr_2_104);

mulc_3_104 : entity work.gfmul
port map(
a=>a_3,
b=>"1100100100",
X=>mulr_3_104);

mulc_4_104 : entity work.gfmul
port map(
a=>a_4,
b=>"0100010000",
X=>mulr_4_104);

mulr_1_105<=a_1;
mulc_2_105 : entity work.gfmul
port map(
a=>a_2,
b=>"1010110000",
X=>mulr_2_105);

mulc_3_105 : entity work.gfmul
port map(
a=>a_3,
b=>"0010001011",
X=>mulr_3_105);

mulc_4_105 : entity work.gfmul
port map(
a=>a_4,
b=>"0010010010",
X=>mulr_4_105);

mulr_1_106<=a_1;
mulc_2_106 : entity work.gfmul
port map(
a=>a_2,
b=>"0101101001",
X=>mulr_2_106);

mulc_3_106 : entity work.gfmul
port map(
a=>a_3,
b=>"1000101100",
X=>mulr_3_106);

mulc_4_106 : entity work.gfmul
port map(
a=>a_4,
b=>"0010011001",
X=>mulr_4_106);

mulr_1_107<=a_1;
mulc_2_107 : entity work.gfmul
port map(
a=>a_2,
b=>"1011010010",
X=>mulr_2_107);

mulc_3_107 : entity work.gfmul
port map(
a=>a_3,
b=>"0010100010",
X=>mulr_3_107);

mulc_4_107 : entity work.gfmul
port map(
a=>a_4,
b=>"0011000001",
X=>mulr_4_107);

mulr_1_108<=a_1;
mulc_2_108 : entity work.gfmul
port map(
a=>a_2,
b=>"0110101101",
X=>mulr_2_108);

mulc_3_108 : entity work.gfmul
port map(
a=>a_3,
b=>"1010001000",
X=>mulr_3_108);

mulc_4_108 : entity work.gfmul
port map(
a=>a_4,
b=>"1000000001",
X=>mulr_4_108);

mulr_1_109<=a_1;
mulc_2_109 : entity work.gfmul
port map(
a=>a_2,
b=>"1101011010",
X=>mulr_2_109);

mulc_3_109 : entity work.gfmul
port map(
a=>a_3,
b=>"1000110010",
X=>mulr_3_109);

mulc_4_109 : entity work.gfmul
port map(
a=>a_4,
b=>"0000101100",
X=>mulr_4_109);

mulr_1_110<=a_1;
mulc_2_110 : entity work.gfmul
port map(
a=>a_2,
b=>"1010111101",
X=>mulr_2_110);

mulc_3_110 : entity work.gfmul
port map(
a=>a_3,
b=>"0011011010",
X=>mulr_3_110);

mulc_4_110 : entity work.gfmul
port map(
a=>a_4,
b=>"0101100000",
X=>mulr_4_110);

mulr_1_111<=a_1;
mulc_2_111 : entity work.gfmul
port map(
a=>a_2,
b=>"0101110011",
X=>mulr_2_111);

mulc_3_111 : entity work.gfmul
port map(
a=>a_3,
b=>"1101101000",
X=>mulr_3_111);

mulc_4_111 : entity work.gfmul
port map(
a=>a_4,
b=>"1100010010",
X=>mulr_4_111);

mulr_1_112<=a_1;
mulc_2_112 : entity work.gfmul
port map(
a=>a_2,
b=>"1011100110",
X=>mulr_2_112);

mulc_3_112 : entity work.gfmul
port map(
a=>a_3,
b=>"0110111011",
X=>mulr_3_112);

mulc_4_112 : entity work.gfmul
port map(
a=>a_4,
b=>"0010100110",
X=>mulr_4_112);

mulr_1_113<=a_1;
mulc_2_113 : entity work.gfmul
port map(
a=>a_2,
b=>"0111000101",
X=>mulr_2_113);

mulc_3_113 : entity work.gfmul
port map(
a=>a_3,
b=>"1011100101",
X=>mulr_3_113);

mulc_4_113 : entity work.gfmul
port map(
a=>a_4,
b=>"0100111001",
X=>mulr_4_113);

mulr_1_114<=a_1;
mulc_2_114 : entity work.gfmul
port map(
a=>a_2,
b=>"1110001010",
X=>mulr_2_114);

mulc_3_114 : entity work.gfmul
port map(
a=>a_3,
b=>"1110000110",
X=>mulr_3_114);

mulc_4_114 : entity work.gfmul
port map(
a=>a_4,
b=>"0111011010",
X=>mulr_4_114);

mulr_1_115<=a_1;
mulc_2_115 : entity work.gfmul
port map(
a=>a_2,
b=>"1100011101",
X=>mulr_2_115);

mulc_3_115 : entity work.gfmul
port map(
a=>a_3,
b=>"1000000011",
X=>mulr_3_115);

mulc_4_115 : entity work.gfmul
port map(
a=>a_4,
b=>"1011001011",
X=>mulr_4_115);

mulr_1_116<=a_1;
mulc_2_116 : entity work.gfmul
port map(
a=>a_2,
b=>"1000110011",
X=>mulr_2_116);

mulc_3_116 : entity work.gfmul
port map(
a=>a_3,
b=>"0000011110",
X=>mulr_3_116);

mulc_4_116 : entity work.gfmul
port map(
a=>a_4,
b=>"1001110101",
X=>mulr_4_116);

mulr_1_117<=a_1;
mulc_2_117 : entity work.gfmul
port map(
a=>a_2,
b=>"0001101111",
X=>mulr_2_117);

mulc_3_117 : entity work.gfmul
port map(
a=>a_3,
b=>"0001111000",
X=>mulr_3_117);

mulc_4_117 : entity work.gfmul
port map(
a=>a_4,
b=>"1110001100",
X=>mulr_4_117);

mulr_1_118<=a_1;
mulc_2_118 : entity work.gfmul
port map(
a=>a_2,
b=>"0011011110",
X=>mulr_2_118);

mulc_3_118 : entity work.gfmul
port map(
a=>a_3,
b=>"0111100000",
X=>mulr_3_118);

mulc_4_118 : entity work.gfmul
port map(
a=>a_4,
b=>"0001011111",
X=>mulr_4_118);

mulr_1_119<=a_1;
mulc_2_119 : entity work.gfmul
port map(
a=>a_2,
b=>"0110111100",
X=>mulr_2_119);

mulc_3_119 : entity work.gfmul
port map(
a=>a_3,
b=>"1110001001",
X=>mulr_3_119);

mulc_4_119 : entity work.gfmul
port map(
a=>a_4,
b=>"1011111000",
X=>mulr_4_119);

mulr_1_120<=a_1;
mulc_2_120 : entity work.gfmul
port map(
a=>a_2,
b=>"1101111000",
X=>mulr_2_120);

mulc_3_120 : entity work.gfmul
port map(
a=>a_3,
b=>"1000111111",
X=>mulr_3_120);

mulc_4_120 : entity work.gfmul
port map(
a=>a_4,
b=>"1111101101",
X=>mulr_4_120);

mulr_1_121<=a_1;
mulc_2_121 : entity work.gfmul
port map(
a=>a_2,
b=>"1011111001",
X=>mulr_2_121);

mulc_3_121 : entity work.gfmul
port map(
a=>a_3,
b=>"0011101110",
X=>mulr_3_121);

mulc_4_121 : entity work.gfmul
port map(
a=>a_4,
b=>"1101010111",
X=>mulr_4_121);

mulr_1_122<=a_1;
mulc_2_122 : entity work.gfmul
port map(
a=>a_2,
b=>"0111111011",
X=>mulr_2_122);

mulc_3_122 : entity work.gfmul
port map(
a=>a_3,
b=>"1110111000",
X=>mulr_3_122);

mulc_4_122 : entity work.gfmul
port map(
a=>a_4,
b=>"1010001110",
X=>mulr_4_122);

mulr_1_123<=a_1;
mulc_2_123 : entity work.gfmul
port map(
a=>a_2,
b=>"1111110110",
X=>mulr_2_123);

mulc_3_123 : entity work.gfmul
port map(
a=>a_3,
b=>"1011111011",
X=>mulr_3_123);

mulc_4_123 : entity work.gfmul
port map(
a=>a_4,
b=>"0001011101",
X=>mulr_4_123);

mulr_1_124<=a_1;
mulc_2_124 : entity work.gfmul
port map(
a=>a_2,
b=>"1111100101",
X=>mulr_2_124);

mulc_3_124 : entity work.gfmul
port map(
a=>a_3,
b=>"1111111110",
X=>mulr_3_124);

mulc_4_124 : entity work.gfmul
port map(
a=>a_4,
b=>"1011101000",
X=>mulr_4_124);

mulr_1_125<=a_1;
mulc_2_125 : entity work.gfmul
port map(
a=>a_2,
b=>"1111000011",
X=>mulr_2_125);

mulc_3_125 : entity work.gfmul
port map(
a=>a_3,
b=>"1111100011",
X=>mulr_3_125);

mulc_4_125 : entity work.gfmul
port map(
a=>a_4,
b=>"1101101101",
X=>mulr_4_125);

mulr_1_126<=a_1;
mulc_2_126 : entity work.gfmul
port map(
a=>a_2,
b=>"1110001111",
X=>mulr_2_126);

mulc_3_126 : entity work.gfmul
port map(
a=>a_3,
b=>"1110010111",
X=>mulr_3_126);

mulc_4_126 : entity work.gfmul
port map(
a=>a_4,
b=>"1101011110",
X=>mulr_4_126);

mulr_1_127<=a_1;
mulc_2_127 : entity work.gfmul
port map(
a=>a_2,
b=>"1100010111",
X=>mulr_2_127);

mulc_3_127 : entity work.gfmul
port map(
a=>a_3,
b=>"1001000111",
X=>mulr_3_127);

mulc_4_127 : entity work.gfmul
port map(
a=>a_4,
b=>"1011000110",
X=>mulr_4_127);

mulr_1_128<=a_1;
mulc_2_128 : entity work.gfmul
port map(
a=>a_2,
b=>"1000100111",
X=>mulr_2_128);

mulc_3_128 : entity work.gfmul
port map(
a=>a_3,
b=>"0100001110",
X=>mulr_3_128);

mulc_4_128 : entity work.gfmul
port map(
a=>a_4,
b=>"1000011101",
X=>mulr_4_128);

mulr_1_129<=a_1;
mulc_2_129 : entity work.gfmul
port map(
a=>a_2,
b=>"0001000111",
X=>mulr_2_129);

mulc_3_129 : entity work.gfmul
port map(
a=>a_3,
b=>"0000110001",
X=>mulr_3_129);

mulc_4_129 : entity work.gfmul
port map(
a=>a_4,
b=>"0011001100",
X=>mulr_4_129);

mulr_1_130<=a_1;
mulc_2_130 : entity work.gfmul
port map(
a=>a_2,
b=>"0010001110",
X=>mulr_2_130);

mulc_3_130 : entity work.gfmul
port map(
a=>a_3,
b=>"0011000100",
X=>mulr_3_130);

mulc_4_130 : entity work.gfmul
port map(
a=>a_4,
b=>"1001101001",
X=>mulr_4_130);

mulr_1_131<=a_1;
mulc_2_131 : entity work.gfmul
port map(
a=>a_2,
b=>"0100011100",
X=>mulr_2_131);

mulc_3_131 : entity work.gfmul
port map(
a=>a_3,
b=>"1100010000",
X=>mulr_3_131);

mulc_4_131 : entity work.gfmul
port map(
a=>a_4,
b=>"1101101100",
X=>mulr_4_131);

mulr_1_132<=a_1;
mulc_2_132 : entity work.gfmul
port map(
a=>a_2,
b=>"1000111000",
X=>mulr_2_132);

mulc_3_132 : entity work.gfmul
port map(
a=>a_3,
b=>"0001011011",
X=>mulr_3_132);

mulc_4_132 : entity work.gfmul
port map(
a=>a_4,
b=>"1101010110",
X=>mulr_4_132);

mulr_1_133<=a_1;
mulc_2_133 : entity work.gfmul
port map(
a=>a_2,
b=>"0001111001",
X=>mulr_2_133);

mulc_3_133 : entity work.gfmul
port map(
a=>a_3,
b=>"0101101100",
X=>mulr_3_133);

mulc_4_133 : entity work.gfmul
port map(
a=>a_4,
b=>"1010000110",
X=>mulr_4_133);

mulr_1_134<=a_1;
mulc_2_134 : entity work.gfmul
port map(
a=>a_2,
b=>"0011110010",
X=>mulr_2_134);

mulc_3_134 : entity work.gfmul
port map(
a=>a_3,
b=>"0110111001",
X=>mulr_3_134);

mulc_4_134 : entity work.gfmul
port map(
a=>a_4,
b=>"0000011101",
X=>mulr_4_134);

mulr_1_135<=a_1;
mulc_2_135 : entity work.gfmul
port map(
a=>a_2,
b=>"0111100100",
X=>mulr_2_135);

mulc_3_135 : entity work.gfmul
port map(
a=>a_3,
b=>"1011101101",
X=>mulr_3_135);

mulc_4_135 : entity work.gfmul
port map(
a=>a_4,
b=>"0011101000",
X=>mulr_4_135);

mulr_1_136<=a_1;
mulc_2_136 : entity work.gfmul
port map(
a=>a_2,
b=>"1111001000",
X=>mulr_2_136);

mulc_3_136 : entity work.gfmul
port map(
a=>a_3,
b=>"1110100110",
X=>mulr_3_136);

mulc_4_136 : entity work.gfmul
port map(
a=>a_4,
b=>"1101001001",
X=>mulr_4_136);

mulr_1_137<=a_1;
mulc_2_137 : entity work.gfmul
port map(
a=>a_2,
b=>"1110011001",
X=>mulr_2_137);

mulc_3_137 : entity work.gfmul
port map(
a=>a_3,
b=>"1010000011",
X=>mulr_3_137);

mulc_4_137 : entity work.gfmul
port map(
a=>a_4,
b=>"1001111110",
X=>mulr_4_137);

mulr_1_138<=a_1;
mulc_2_138 : entity work.gfmul
port map(
a=>a_2,
b=>"1100111011",
X=>mulr_2_138);

mulc_3_138 : entity work.gfmul
port map(
a=>a_3,
b=>"1000011110",
X=>mulr_3_138);

mulc_4_138 : entity work.gfmul
port map(
a=>a_4,
b=>"1111010100",
X=>mulr_4_138);

mulr_1_139<=a_1;
mulc_2_139 : entity work.gfmul
port map(
a=>a_2,
b=>"1001111111",
X=>mulr_2_139);

mulc_3_139 : entity work.gfmul
port map(
a=>a_3,
b=>"0001101010",
X=>mulr_3_139);

mulc_4_139 : entity work.gfmul
port map(
a=>a_4,
b=>"1010011111",
X=>mulr_4_139);

mulr_1_140<=a_1;
mulc_2_140 : entity work.gfmul
port map(
a=>a_2,
b=>"0011110111",
X=>mulr_2_140);

mulc_3_140 : entity work.gfmul
port map(
a=>a_3,
b=>"0110101000",
X=>mulr_3_140);

mulc_4_140 : entity work.gfmul
port map(
a=>a_4,
b=>"0011010101",
X=>mulr_4_140);

mulr_1_141<=a_1;
mulc_2_141 : entity work.gfmul
port map(
a=>a_2,
b=>"0111101110",
X=>mulr_2_141);

mulc_3_141 : entity work.gfmul
port map(
a=>a_3,
b=>"1010101001",
X=>mulr_3_141);

mulc_4_141 : entity work.gfmul
port map(
a=>a_4,
b=>"1010100001",
X=>mulr_4_141);

mulr_1_142<=a_1;
mulc_2_142 : entity work.gfmul
port map(
a=>a_2,
b=>"1111011100",
X=>mulr_2_142);

mulc_3_142 : entity work.gfmul
port map(
a=>a_3,
b=>"1010110110",
X=>mulr_3_142);

mulc_4_142 : entity work.gfmul
port map(
a=>a_4,
b=>"0100100101",
X=>mulr_4_142);

mulr_1_143<=a_1;
mulc_2_143 : entity work.gfmul
port map(
a=>a_2,
b=>"1110110001",
X=>mulr_2_143);

mulc_3_143 : entity work.gfmul
port map(
a=>a_3,
b=>"1011001010",
X=>mulr_3_143);

mulc_4_143 : entity work.gfmul
port map(
a=>a_4,
b=>"0100111010",
X=>mulr_4_143);

mulr_1_144<=a_1;
mulc_2_144 : entity work.gfmul
port map(
a=>a_2,
b=>"1101101011",
X=>mulr_2_144);

mulc_3_144 : entity work.gfmul
port map(
a=>a_3,
b=>"1100111010",
X=>mulr_3_144);

mulc_4_144 : entity work.gfmul
port map(
a=>a_4,
b=>"0111000010",
X=>mulr_4_144);

mulr_1_145<=a_1;
mulc_2_145 : entity work.gfmul
port map(
a=>a_2,
b=>"1011011111",
X=>mulr_2_145);

mulc_3_145 : entity work.gfmul
port map(
a=>a_3,
b=>"0011110011",
X=>mulr_3_145);

mulc_4_145 : entity work.gfmul
port map(
a=>a_4,
b=>"1000001011",
X=>mulr_4_145);

mulr_1_146<=a_1;
mulc_2_146 : entity work.gfmul
port map(
a=>a_2,
b=>"0110110111",
X=>mulr_2_146);

mulc_3_146 : entity work.gfmul
port map(
a=>a_3,
b=>"1111001100",
X=>mulr_3_146);

mulc_4_146 : entity work.gfmul
port map(
a=>a_4,
b=>"0001111100",
X=>mulr_4_146);

mulr_1_147<=a_1;
mulc_2_147 : entity work.gfmul
port map(
a=>a_2,
b=>"1101101110",
X=>mulr_2_147);

mulc_3_147 : entity work.gfmul
port map(
a=>a_3,
b=>"1100101011",
X=>mulr_3_147);

mulc_4_147 : entity work.gfmul
port map(
a=>a_4,
b=>"1111100000",
X=>mulr_4_147);

mulr_1_148<=a_1;
mulc_2_148 : entity work.gfmul
port map(
a=>a_2,
b=>"1011010101",
X=>mulr_2_148);

mulc_3_148 : entity work.gfmul
port map(
a=>a_3,
b=>"0010110111",
X=>mulr_3_148);

mulc_4_148 : entity work.gfmul
port map(
a=>a_4,
b=>"1100111111",
X=>mulr_4_148);

mulr_1_149<=a_1;
mulc_2_149 : entity work.gfmul
port map(
a=>a_2,
b=>"0110100011",
X=>mulr_2_149);

mulc_3_149 : entity work.gfmul
port map(
a=>a_3,
b=>"1011011100",
X=>mulr_3_149);

mulc_4_149 : entity work.gfmul
port map(
a=>a_4,
b=>"0111001110",
X=>mulr_4_149);

mulr_1_150<=a_1;
mulc_2_150 : entity work.gfmul
port map(
a=>a_2,
b=>"1101000110",
X=>mulr_2_150);

mulc_3_150 : entity work.gfmul
port map(
a=>a_3,
b=>"1101100010",
X=>mulr_3_150);

mulc_4_150 : entity work.gfmul
port map(
a=>a_4,
b=>"1001101011",
X=>mulr_4_150);

mulr_1_151<=a_1;
mulc_2_151 : entity work.gfmul
port map(
a=>a_2,
b=>"1010000101",
X=>mulr_2_151);

mulc_3_151 : entity work.gfmul
port map(
a=>a_3,
b=>"0110010011",
X=>mulr_3_151);

mulc_4_151 : entity work.gfmul
port map(
a=>a_4,
b=>"1101111100",
X=>mulr_4_151);

mulr_1_152<=a_1;
mulc_2_152 : entity work.gfmul
port map(
a=>a_2,
b=>"0100000011",
X=>mulr_2_152);

mulc_3_152 : entity work.gfmul
port map(
a=>a_3,
b=>"1001000101",
X=>mulr_3_152);

mulc_4_152 : entity work.gfmul
port map(
a=>a_4,
b=>"1111010110",
X=>mulr_4_152);

mulr_1_153<=a_1;
mulc_2_153 : entity work.gfmul
port map(
a=>a_2,
b=>"1000000110",
X=>mulr_2_153);

mulc_3_153 : entity work.gfmul
port map(
a=>a_3,
b=>"0100000110",
X=>mulr_3_153);

mulc_4_153 : entity work.gfmul
port map(
a=>a_4,
b=>"1010001111",
X=>mulr_4_153);

mulr_1_154<=a_1;
mulc_2_154 : entity work.gfmul
port map(
a=>a_2,
b=>"0000000101",
X=>mulr_2_154);

mulc_3_154 : entity work.gfmul
port map(
a=>a_3,
b=>"0000010001",
X=>mulr_3_154);

mulc_4_154 : entity work.gfmul
port map(
a=>a_4,
b=>"0001010101",
X=>mulr_4_154);

mulr_1_155<=a_1;
mulc_2_155 : entity work.gfmul
port map(
a=>a_2,
b=>"0000001010",
X=>mulr_2_155);

mulc_3_155 : entity work.gfmul
port map(
a=>a_3,
b=>"0001000100",
X=>mulr_3_155);

mulc_4_155 : entity work.gfmul
port map(
a=>a_4,
b=>"1010101000",
X=>mulr_4_155);

mulr_1_156<=a_1;
mulc_2_156 : entity work.gfmul
port map(
a=>a_2,
b=>"0000010100",
X=>mulr_2_156);

mulc_3_156 : entity work.gfmul
port map(
a=>a_3,
b=>"0100010000",
X=>mulr_3_156);

mulc_4_156 : entity work.gfmul
port map(
a=>a_4,
b=>"0101101101",
X=>mulr_4_156);

mulr_1_157<=a_1;
mulc_2_157 : entity work.gfmul
port map(
a=>a_2,
b=>"0000101000",
X=>mulr_2_157);

mulc_3_157 : entity work.gfmul
port map(
a=>a_3,
b=>"0001001001",
X=>mulr_3_157);

mulc_4_157 : entity work.gfmul
port map(
a=>a_4,
b=>"1101111010",
X=>mulr_4_157);

mulr_1_158<=a_1;
mulc_2_158 : entity work.gfmul
port map(
a=>a_2,
b=>"0001010000",
X=>mulr_2_158);

mulc_3_158 : entity work.gfmul
port map(
a=>a_3,
b=>"0100100100",
X=>mulr_3_158);

mulc_4_158 : entity work.gfmul
port map(
a=>a_4,
b=>"1111100110",
X=>mulr_4_158);

mulr_1_159<=a_1;
mulc_2_159 : entity work.gfmul
port map(
a=>a_2,
b=>"0010100000",
X=>mulr_2_159);

mulc_3_159 : entity work.gfmul
port map(
a=>a_3,
b=>"0010011001",
X=>mulr_3_159);

mulc_4_159 : entity work.gfmul
port map(
a=>a_4,
b=>"1100001111",
X=>mulr_4_159);

mulr_1_160<=a_1;
mulc_2_160 : entity work.gfmul
port map(
a=>a_2,
b=>"0101000000",
X=>mulr_2_160);

mulc_3_160 : entity work.gfmul
port map(
a=>a_3,
b=>"1001100100",
X=>mulr_3_160);

mulc_4_160 : entity work.gfmul
port map(
a=>a_4,
b=>"0001001110",
X=>mulr_4_160);

mulr_1_161<=a_1;
mulc_2_161 : entity work.gfmul
port map(
a=>a_2,
b=>"1010000000",
X=>mulr_2_161);

mulc_3_161 : entity work.gfmul
port map(
a=>a_3,
b=>"0110000010",
X=>mulr_3_161);

mulc_4_161 : entity work.gfmul
port map(
a=>a_4,
b=>"1001110000",
X=>mulr_4_161);

mulr_1_162<=a_1;
mulc_2_162 : entity work.gfmul
port map(
a=>a_2,
b=>"0100001001",
X=>mulr_2_162);

mulc_3_162 : entity work.gfmul
port map(
a=>a_3,
b=>"1000000001",
X=>mulr_3_162);

mulc_4_162 : entity work.gfmul
port map(
a=>a_4,
b=>"1110100100",
X=>mulr_4_162);

mulr_1_163<=a_1;
mulc_2_163 : entity work.gfmul
port map(
a=>a_2,
b=>"1000010010",
X=>mulr_2_163);

mulc_3_163 : entity work.gfmul
port map(
a=>a_3,
b=>"0000010110",
X=>mulr_3_163);

mulc_4_163 : entity work.gfmul
port map(
a=>a_4,
b=>"0100011111",
X=>mulr_4_163);

mulr_1_164<=a_1;
mulc_2_164 : entity work.gfmul
port map(
a=>a_2,
b=>"0000101101",
X=>mulr_2_164);

mulc_3_164 : entity work.gfmul
port map(
a=>a_3,
b=>"0001011000",
X=>mulr_3_164);

mulc_4_164 : entity work.gfmul
port map(
a=>a_4,
b=>"0011101010",
X=>mulr_4_164);

mulr_1_165<=a_1;
mulc_2_165 : entity work.gfmul
port map(
a=>a_2,
b=>"0001011010",
X=>mulr_2_165);

mulc_3_165 : entity work.gfmul
port map(
a=>a_3,
b=>"0101100000",
X=>mulr_3_165);

mulc_4_165 : entity work.gfmul
port map(
a=>a_4,
b=>"1101011001",
X=>mulr_4_165);

mulr_1_166<=a_1;
mulc_2_166 : entity work.gfmul
port map(
a=>a_2,
b=>"0010110100",
X=>mulr_2_166);

mulc_3_166 : entity work.gfmul
port map(
a=>a_3,
b=>"0110001001",
X=>mulr_3_166);

mulc_4_166 : entity work.gfmul
port map(
a=>a_4,
b=>"1011111110",
X=>mulr_4_166);

mulr_1_167<=a_1;
mulc_2_167 : entity work.gfmul
port map(
a=>a_2,
b=>"0101101000",
X=>mulr_2_167);

mulc_3_167 : entity work.gfmul
port map(
a=>a_3,
b=>"1000101101",
X=>mulr_3_167);

mulc_4_167 : entity work.gfmul
port map(
a=>a_4,
b=>"1111011101",
X=>mulr_4_167);

mulr_1_168<=a_1;
mulc_2_168 : entity work.gfmul
port map(
a=>a_2,
b=>"1011010000",
X=>mulr_2_168);

mulc_3_168 : entity work.gfmul
port map(
a=>a_3,
b=>"0010100110",
X=>mulr_3_168);

mulc_4_168 : entity work.gfmul
port map(
a=>a_4,
b=>"1011010111",
X=>mulr_4_168);

mulr_1_169<=a_1;
mulc_2_169 : entity work.gfmul
port map(
a=>a_2,
b=>"0110101001",
X=>mulr_2_169);

mulc_3_169 : entity work.gfmul
port map(
a=>a_3,
b=>"1010011000",
X=>mulr_3_169);

mulc_4_169 : entity work.gfmul
port map(
a=>a_4,
b=>"1010010101",
X=>mulr_4_169);

mulr_1_170<=a_1;
mulc_2_170 : entity work.gfmul
port map(
a=>a_2,
b=>"1101010010",
X=>mulr_2_170);

mulc_3_170 : entity work.gfmul
port map(
a=>a_3,
b=>"1001110010",
X=>mulr_3_170);

mulc_4_170 : entity work.gfmul
port map(
a=>a_4,
b=>"0010000101",
X=>mulr_4_170);

mulr_1_171<=a_1;
mulc_2_171 : entity work.gfmul
port map(
a=>a_2,
b=>"1010101101",
X=>mulr_2_171);

mulc_3_171 : entity work.gfmul
port map(
a=>a_3,
b=>"0111011010",
X=>mulr_3_171);

mulc_4_171 : entity work.gfmul
port map(
a=>a_4,
b=>"0000100001",
X=>mulr_4_171);

mulr_1_172<=a_1;
mulc_2_172 : entity work.gfmul
port map(
a=>a_2,
b=>"0101010011",
X=>mulr_2_172);

mulc_3_172 : entity work.gfmul
port map(
a=>a_3,
b=>"1101100001",
X=>mulr_3_172);

mulc_4_172 : entity work.gfmul
port map(
a=>a_4,
b=>"0100001000",
X=>mulr_4_172);

mulr_1_173<=a_1;
mulc_2_173 : entity work.gfmul
port map(
a=>a_2,
b=>"1010100110",
X=>mulr_2_173);

mulc_3_173 : entity work.gfmul
port map(
a=>a_3,
b=>"0110011111",
X=>mulr_3_173);

mulc_4_173 : entity work.gfmul
port map(
a=>a_4,
b=>"0001010010",
X=>mulr_4_173);

mulr_1_174<=a_1;
mulc_2_174 : entity work.gfmul
port map(
a=>a_2,
b=>"0101000101",
X=>mulr_2_174);

mulc_3_174 : entity work.gfmul
port map(
a=>a_3,
b=>"1001110101",
X=>mulr_3_174);

mulc_4_174 : entity work.gfmul
port map(
a=>a_4,
b=>"1010010000",
X=>mulr_4_174);

mulr_1_175<=a_1;
mulc_2_175 : entity work.gfmul
port map(
a=>a_2,
b=>"1010001010",
X=>mulr_2_175);

mulc_3_175 : entity work.gfmul
port map(
a=>a_3,
b=>"0111000110",
X=>mulr_3_175);

mulc_4_175 : entity work.gfmul
port map(
a=>a_4,
b=>"0010101101",
X=>mulr_4_175);

mulr_1_176<=a_1;
mulc_2_176 : entity work.gfmul
port map(
a=>a_2,
b=>"0100011101",
X=>mulr_2_176);

mulc_3_176 : entity work.gfmul
port map(
a=>a_3,
b=>"1100010001",
X=>mulr_3_176);

mulc_4_176 : entity work.gfmul
port map(
a=>a_4,
b=>"0101100001",
X=>mulr_4_176);

mulr_1_177<=a_1;
mulc_2_177 : entity work.gfmul
port map(
a=>a_2,
b=>"1000111010",
X=>mulr_2_177);

mulc_3_177 : entity work.gfmul
port map(
a=>a_3,
b=>"0001011111",
X=>mulr_3_177);

mulc_4_177 : entity work.gfmul
port map(
a=>a_4,
b=>"1100011010",
X=>mulr_4_177);

mulr_1_178<=a_1;
mulc_2_178 : entity work.gfmul
port map(
a=>a_2,
b=>"0001111101",
X=>mulr_2_178);

mulc_3_178 : entity work.gfmul
port map(
a=>a_3,
b=>"0101111100",
X=>mulr_3_178);

mulc_4_178 : entity work.gfmul
port map(
a=>a_4,
b=>"0011100110",
X=>mulr_4_178);

mulr_1_179<=a_1;
mulc_2_179 : entity work.gfmul
port map(
a=>a_2,
b=>"0011111010",
X=>mulr_2_179);

mulc_3_179 : entity work.gfmul
port map(
a=>a_3,
b=>"0111111001",
X=>mulr_3_179);

mulc_4_179 : entity work.gfmul
port map(
a=>a_4,
b=>"1100111001",
X=>mulr_4_179);

mulr_1_180<=a_1;
mulc_2_180 : entity work.gfmul
port map(
a=>a_2,
b=>"0111110100",
X=>mulr_2_180);

mulc_3_180 : entity work.gfmul
port map(
a=>a_3,
b=>"1111101101",
X=>mulr_3_180);

mulc_4_180 : entity work.gfmul
port map(
a=>a_4,
b=>"0111111110",
X=>mulr_4_180);

mulr_1_181<=a_1;
mulc_2_181 : entity work.gfmul
port map(
a=>a_2,
b=>"1111101000",
X=>mulr_2_181);

mulc_3_181 : entity work.gfmul
port map(
a=>a_3,
b=>"1110101111",
X=>mulr_3_181);

mulc_4_181 : entity work.gfmul
port map(
a=>a_4,
b=>"1111101011",
X=>mulr_4_181);

mulr_1_182<=a_1;
mulc_2_182 : entity work.gfmul
port map(
a=>a_2,
b=>"1111011001",
X=>mulr_2_182);

mulc_3_182 : entity work.gfmul
port map(
a=>a_3,
b=>"1010100111",
X=>mulr_3_182);

mulc_4_182 : entity work.gfmul
port map(
a=>a_4,
b=>"1101100111",
X=>mulr_4_182);

mulr_1_183<=a_1;
mulc_2_183 : entity work.gfmul
port map(
a=>a_2,
b=>"1110111011",
X=>mulr_2_183);

mulc_3_183 : entity work.gfmul
port map(
a=>a_3,
b=>"1010001110",
X=>mulr_3_183);

mulc_4_183 : entity work.gfmul
port map(
a=>a_4,
b=>"1100001110",
X=>mulr_4_183);

mulr_1_184<=a_1;
mulc_2_184 : entity work.gfmul
port map(
a=>a_2,
b=>"1101111111",
X=>mulr_2_184);

mulc_3_184 : entity work.gfmul
port map(
a=>a_3,
b=>"1000101010",
X=>mulr_3_184);

mulc_4_184 : entity work.gfmul
port map(
a=>a_4,
b=>"0001000110",
X=>mulr_4_184);

mulr_1_185<=a_1;
mulc_2_185 : entity work.gfmul
port map(
a=>a_2,
b=>"1011110111",
X=>mulr_2_185);

mulc_3_185 : entity work.gfmul
port map(
a=>a_3,
b=>"0010111010",
X=>mulr_3_185);

mulc_4_185 : entity work.gfmul
port map(
a=>a_4,
b=>"1000110000",
X=>mulr_4_185);

mulr_1_186<=a_1;
mulc_2_186 : entity work.gfmul
port map(
a=>a_2,
b=>"0111100111",
X=>mulr_2_186);

mulc_3_186 : entity work.gfmul
port map(
a=>a_3,
b=>"1011101000",
X=>mulr_3_186);

mulc_4_186 : entity work.gfmul
port map(
a=>a_4,
b=>"0110100100",
X=>mulr_4_186);

mulr_1_187<=a_1;
mulc_2_187 : entity work.gfmul
port map(
a=>a_2,
b=>"1111001110",
X=>mulr_2_187);

mulc_3_187 : entity work.gfmul
port map(
a=>a_3,
b=>"1110110010",
X=>mulr_3_187);

mulc_4_187 : entity work.gfmul
port map(
a=>a_4,
b=>"0100111011",
X=>mulr_4_187);

mulr_1_188<=a_1;
mulc_2_188 : entity work.gfmul
port map(
a=>a_2,
b=>"1110010101",
X=>mulr_2_188);

mulc_3_188 : entity work.gfmul
port map(
a=>a_3,
b=>"1011010011",
X=>mulr_3_188);

mulc_4_188 : entity work.gfmul
port map(
a=>a_4,
b=>"0111001010",
X=>mulr_4_188);

mulr_1_189<=a_1;
mulc_2_189 : entity work.gfmul
port map(
a=>a_2,
b=>"1100100011",
X=>mulr_2_189);

mulc_3_189 : entity work.gfmul
port map(
a=>a_3,
b=>"1101011110",
X=>mulr_3_189);

mulc_4_189 : entity work.gfmul
port map(
a=>a_4,
b=>"1001001011",
X=>mulr_4_189);

mulr_1_190<=a_1;
mulc_2_190 : entity work.gfmul
port map(
a=>a_2,
b=>"1001001111",
X=>mulr_2_190);

mulc_3_190 : entity work.gfmul
port map(
a=>a_3,
b=>"0101100011",
X=>mulr_3_190);

mulc_4_190 : entity work.gfmul
port map(
a=>a_4,
b=>"1001111100",
X=>mulr_4_190);

mulr_1_191<=a_1;
mulc_2_191 : entity work.gfmul
port map(
a=>a_2,
b=>"0010010111",
X=>mulr_2_191);

mulc_3_191 : entity work.gfmul
port map(
a=>a_3,
b=>"0110000101",
X=>mulr_3_191);

mulc_4_191 : entity work.gfmul
port map(
a=>a_4,
b=>"1111000100",
X=>mulr_4_191);

mulr_1_192<=a_1;
mulc_2_192 : entity work.gfmul
port map(
a=>a_2,
b=>"0100101110",
X=>mulr_2_192);

mulc_3_192 : entity work.gfmul
port map(
a=>a_3,
b=>"1000011101",
X=>mulr_3_192);

mulc_4_192 : entity work.gfmul
port map(
a=>a_4,
b=>"1000011111",
X=>mulr_4_192);

mulr_1_193<=a_1;
mulc_2_193 : entity work.gfmul
port map(
a=>a_2,
b=>"1001011100",
X=>mulr_2_193);

mulc_3_193 : entity work.gfmul
port map(
a=>a_3,
b=>"0001100110",
X=>mulr_3_193);

mulc_4_193 : entity work.gfmul
port map(
a=>a_4,
b=>"0011011100",
X=>mulr_4_193);

mulr_1_194<=a_1;
mulc_2_194 : entity work.gfmul
port map(
a=>a_2,
b=>"0010110001",
X=>mulr_2_194);

mulc_3_194 : entity work.gfmul
port map(
a=>a_3,
b=>"0110011000",
X=>mulr_3_194);

mulc_4_194 : entity work.gfmul
port map(
a=>a_4,
b=>"1011101001",
X=>mulr_4_194);

mulr_1_195<=a_1;
mulc_2_195 : entity work.gfmul
port map(
a=>a_2,
b=>"0101100010",
X=>mulr_2_195);

mulc_3_195 : entity work.gfmul
port map(
a=>a_3,
b=>"1001101001",
X=>mulr_3_195);

mulc_4_195 : entity work.gfmul
port map(
a=>a_4,
b=>"1101100101",
X=>mulr_4_195);

mulr_1_196<=a_1;
mulc_2_196 : entity work.gfmul
port map(
a=>a_2,
b=>"1011000100",
X=>mulr_2_196);

mulc_3_196 : entity work.gfmul
port map(
a=>a_3,
b=>"0110110110",
X=>mulr_3_196);

mulc_4_196 : entity work.gfmul
port map(
a=>a_4,
b=>"1100011110",
X=>mulr_4_196);

mulr_1_197<=a_1;
mulc_2_197 : entity work.gfmul
port map(
a=>a_2,
b=>"0110000001",
X=>mulr_2_197);

mulc_3_197 : entity work.gfmul
port map(
a=>a_3,
b=>"1011010001",
X=>mulr_3_197);

mulc_4_197 : entity work.gfmul
port map(
a=>a_4,
b=>"0011000110",
X=>mulr_4_197);

mulr_1_198<=a_1;
mulc_2_198 : entity work.gfmul
port map(
a=>a_2,
b=>"1100000010",
X=>mulr_2_198);

mulc_3_198 : entity work.gfmul
port map(
a=>a_3,
b=>"1101010110",
X=>mulr_3_198);

mulc_4_198 : entity work.gfmul
port map(
a=>a_4,
b=>"1000111001",
X=>mulr_4_198);

mulr_1_199<=a_1;
mulc_2_199 : entity work.gfmul
port map(
a=>a_2,
b=>"1000001101",
X=>mulr_2_199);

mulc_3_199 : entity work.gfmul
port map(
a=>a_3,
b=>"0101000011",
X=>mulr_3_199);

mulc_4_199 : entity work.gfmul
port map(
a=>a_4,
b=>"0111101100",
X=>mulr_4_199);

mulr_1_200<=a_1;
mulc_2_200 : entity work.gfmul
port map(
a=>a_2,
b=>"0000010011",
X=>mulr_2_200);

mulc_3_200 : entity work.gfmul
port map(
a=>a_3,
b=>"0100000101",
X=>mulr_3_200);

mulc_4_200 : entity work.gfmul
port map(
a=>a_4,
b=>"1101111011",
X=>mulr_4_200);

mulr_1_201<=a_1;
mulc_2_201 : entity work.gfmul
port map(
a=>a_2,
b=>"0000100110",
X=>mulr_2_201);

mulc_3_201 : entity work.gfmul
port map(
a=>a_3,
b=>"0000011101",
X=>mulr_3_201);

mulc_4_201 : entity work.gfmul
port map(
a=>a_4,
b=>"1111101110",
X=>mulr_4_201);

mulr_1_202<=a_1;
mulc_2_202 : entity work.gfmul
port map(
a=>a_2,
b=>"0001001100",
X=>mulr_2_202);

mulc_3_202 : entity work.gfmul
port map(
a=>a_3,
b=>"0001110100",
X=>mulr_3_202);

mulc_4_202 : entity work.gfmul
port map(
a=>a_4,
b=>"1101001111",
X=>mulr_4_202);

mulr_1_203<=a_1;
mulc_2_203 : entity work.gfmul
port map(
a=>a_2,
b=>"0010011000",
X=>mulr_2_203);

mulc_3_203 : entity work.gfmul
port map(
a=>a_3,
b=>"0111010000",
X=>mulr_3_203);

mulc_4_203 : entity work.gfmul
port map(
a=>a_4,
b=>"1001001110",
X=>mulr_4_203);

mulr_1_204<=a_1;
mulc_2_204 : entity work.gfmul
port map(
a=>a_2,
b=>"0100110000",
X=>mulr_2_204);

mulc_3_204 : entity work.gfmul
port map(
a=>a_3,
b=>"1101001001",
X=>mulr_3_204);

mulc_4_204 : entity work.gfmul
port map(
a=>a_4,
b=>"1001010100",
X=>mulr_4_204);

mulr_1_205<=a_1;
mulc_2_205 : entity work.gfmul
port map(
a=>a_2,
b=>"1001100000",
X=>mulr_2_205);

mulc_3_205 : entity work.gfmul
port map(
a=>a_3,
b=>"0100111111",
X=>mulr_3_205);

mulc_4_205 : entity work.gfmul
port map(
a=>a_4,
b=>"1010000100",
X=>mulr_4_205);

mulr_1_206<=a_1;
mulc_2_206 : entity work.gfmul
port map(
a=>a_2,
b=>"0011001001",
X=>mulr_2_206);

mulc_3_206 : entity work.gfmul
port map(
a=>a_3,
b=>"0011110101",
X=>mulr_3_206);

mulc_4_206 : entity work.gfmul
port map(
a=>a_4,
b=>"0000001101",
X=>mulr_4_206);

mulr_1_207<=a_1;
mulc_2_207 : entity work.gfmul
port map(
a=>a_2,
b=>"0110010010",
X=>mulr_2_207);

mulc_3_207 : entity work.gfmul
port map(
a=>a_3,
b=>"1111010100",
X=>mulr_3_207);

mulc_4_207 : entity work.gfmul
port map(
a=>a_4,
b=>"0001101000",
X=>mulr_4_207);

mulr_1_208<=a_1;
mulc_2_208 : entity work.gfmul
port map(
a=>a_2,
b=>"1100100100",
X=>mulr_2_208);

mulc_3_208 : entity work.gfmul
port map(
a=>a_3,
b=>"1101001011",
X=>mulr_3_208);

mulc_4_208 : entity work.gfmul
port map(
a=>a_4,
b=>"1101000000",
X=>mulr_4_208);

mulr_1_209<=a_1;
mulc_2_209 : entity work.gfmul
port map(
a=>a_2,
b=>"1001000001",
X=>mulr_2_209);

mulc_3_209 : entity work.gfmul
port map(
a=>a_3,
b=>"0100110111",
X=>mulr_3_209);

mulc_4_209 : entity work.gfmul
port map(
a=>a_4,
b=>"1000110110",
X=>mulr_4_209);

mulr_1_210<=a_1;
mulc_2_210 : entity work.gfmul
port map(
a=>a_2,
b=>"0010001011",
X=>mulr_2_210);

mulc_3_210 : entity work.gfmul
port map(
a=>a_3,
b=>"0011010101",
X=>mulr_3_210);

mulc_4_210 : entity work.gfmul
port map(
a=>a_4,
b=>"0110010100",
X=>mulr_4_210);

mulr_1_211<=a_1;
mulc_2_211 : entity work.gfmul
port map(
a=>a_2,
b=>"0100010110",
X=>mulr_2_211);

mulc_3_211 : entity work.gfmul
port map(
a=>a_3,
b=>"1101010100",
X=>mulr_3_211);

mulc_4_211 : entity work.gfmul
port map(
a=>a_4,
b=>"0010111011",
X=>mulr_4_211);

mulr_1_212<=a_1;
mulc_2_212 : entity work.gfmul
port map(
a=>a_2,
b=>"1000101100",
X=>mulr_2_212);

mulc_3_212 : entity work.gfmul
port map(
a=>a_3,
b=>"0101001011",
X=>mulr_3_212);

mulc_4_212 : entity work.gfmul
port map(
a=>a_4,
b=>"0111010001",
X=>mulr_4_212);

mulr_1_213<=a_1;
mulc_2_213 : entity work.gfmul
port map(
a=>a_2,
b=>"0001010001",
X=>mulr_2_213);

mulc_3_213 : entity work.gfmul
port map(
a=>a_3,
b=>"0100100101",
X=>mulr_3_213);

mulc_4_213 : entity work.gfmul
port map(
a=>a_4,
b=>"1010010011",
X=>mulr_4_213);

mulr_1_214<=a_1;
mulc_2_214 : entity work.gfmul
port map(
a=>a_2,
b=>"0010100010",
X=>mulr_2_214);

mulc_3_214 : entity work.gfmul
port map(
a=>a_3,
b=>"0010011101",
X=>mulr_3_214);

mulc_4_214 : entity work.gfmul
port map(
a=>a_4,
b=>"0010110101",
X=>mulr_4_214);

mulr_1_215<=a_1;
mulc_2_215 : entity work.gfmul
port map(
a=>a_2,
b=>"0101000100",
X=>mulr_2_215);

mulc_3_215 : entity work.gfmul
port map(
a=>a_3,
b=>"1001110100",
X=>mulr_3_215);

mulc_4_215 : entity work.gfmul
port map(
a=>a_4,
b=>"0110100001",
X=>mulr_4_215);

mulr_1_216<=a_1;
mulc_2_216 : entity work.gfmul
port map(
a=>a_2,
b=>"1010001000",
X=>mulr_2_216);

mulc_3_216 : entity work.gfmul
port map(
a=>a_3,
b=>"0111000010",
X=>mulr_3_216);

mulc_4_216 : entity work.gfmul
port map(
a=>a_4,
b=>"0100010011",
X=>mulr_4_216);

mulr_1_217<=a_1;
mulc_2_217 : entity work.gfmul
port map(
a=>a_2,
b=>"0100011001",
X=>mulr_2_217);

mulc_3_217 : entity work.gfmul
port map(
a=>a_3,
b=>"1100000001",
X=>mulr_3_217);

mulc_4_217 : entity work.gfmul
port map(
a=>a_4,
b=>"0010001010",
X=>mulr_4_217);

mulr_1_218<=a_1;
mulc_2_218 : entity work.gfmul
port map(
a=>a_2,
b=>"1000110010",
X=>mulr_2_218);

mulc_3_218 : entity work.gfmul
port map(
a=>a_3,
b=>"0000011111",
X=>mulr_3_218);

mulc_4_218 : entity work.gfmul
port map(
a=>a_4,
b=>"0001011001",
X=>mulr_4_218);

mulr_1_219<=a_1;
mulc_2_219 : entity work.gfmul
port map(
a=>a_2,
b=>"0001101101",
X=>mulr_2_219);

mulc_3_219 : entity work.gfmul
port map(
a=>a_3,
b=>"0001111100",
X=>mulr_3_219);

mulc_4_219 : entity work.gfmul
port map(
a=>a_4,
b=>"1011001000",
X=>mulr_4_219);

mulr_1_220<=a_1;
mulc_2_220 : entity work.gfmul
port map(
a=>a_2,
b=>"0011011010",
X=>mulr_2_220);

mulc_3_220 : entity work.gfmul
port map(
a=>a_3,
b=>"0111110000",
X=>mulr_3_220);

mulc_4_220 : entity work.gfmul
port map(
a=>a_4,
b=>"1001101101",
X=>mulr_4_220);

mulr_1_221<=a_1;
mulc_2_221 : entity work.gfmul
port map(
a=>a_2,
b=>"0110110100",
X=>mulr_2_221);

mulc_3_221 : entity work.gfmul
port map(
a=>a_3,
b=>"1111001001",
X=>mulr_3_221);

mulc_4_221 : entity work.gfmul
port map(
a=>a_4,
b=>"1101001100",
X=>mulr_4_221);

mulr_1_222<=a_1;
mulc_2_222 : entity work.gfmul
port map(
a=>a_2,
b=>"1101101000",
X=>mulr_2_222);

mulc_3_222 : entity work.gfmul
port map(
a=>a_3,
b=>"1100111111",
X=>mulr_3_222);

mulc_4_222 : entity work.gfmul
port map(
a=>a_4,
b=>"1001010110",
X=>mulr_4_222);

mulr_1_223<=a_1;
mulc_2_223 : entity work.gfmul
port map(
a=>a_2,
b=>"1011011001",
X=>mulr_2_223);

mulc_3_223 : entity work.gfmul
port map(
a=>a_3,
b=>"0011100111",
X=>mulr_3_223);

mulc_4_223 : entity work.gfmul
port map(
a=>a_4,
b=>"1010010100",
X=>mulr_4_223);

mulr_1_224<=a_1;
mulc_2_224 : entity work.gfmul
port map(
a=>a_2,
b=>"0110111011",
X=>mulr_2_224);

mulc_3_224 : entity work.gfmul
port map(
a=>a_3,
b=>"1110011100",
X=>mulr_3_224);

mulc_4_224 : entity work.gfmul
port map(
a=>a_4,
b=>"0010001101",
X=>mulr_4_224);

mulr_1_225<=a_1;
mulc_2_225 : entity work.gfmul
port map(
a=>a_2,
b=>"1101110110",
X=>mulr_2_225);

mulc_3_225 : entity work.gfmul
port map(
a=>a_3,
b=>"1001101011",
X=>mulr_3_225);

mulc_4_225 : entity work.gfmul
port map(
a=>a_4,
b=>"0001100001",
X=>mulr_4_225);

mulr_1_226<=a_1;
mulc_2_226 : entity work.gfmul
port map(
a=>a_2,
b=>"1011100101",
X=>mulr_2_226);

mulc_3_226 : entity work.gfmul
port map(
a=>a_3,
b=>"0110111110",
X=>mulr_3_226);

mulc_4_226 : entity work.gfmul
port map(
a=>a_4,
b=>"1100001000",
X=>mulr_4_226);

mulr_1_227<=a_1;
mulc_2_227 : entity work.gfmul
port map(
a=>a_2,
b=>"0111000011",
X=>mulr_2_227);

mulc_3_227 : entity work.gfmul
port map(
a=>a_3,
b=>"1011110001",
X=>mulr_3_227);

mulc_4_227 : entity work.gfmul
port map(
a=>a_4,
b=>"0001110110",
X=>mulr_4_227);

mulr_1_228<=a_1;
mulc_2_228 : entity work.gfmul
port map(
a=>a_2,
b=>"1110000110",
X=>mulr_2_228);

mulc_3_228 : entity work.gfmul
port map(
a=>a_3,
b=>"1111010110",
X=>mulr_3_228);

mulc_4_228 : entity work.gfmul
port map(
a=>a_4,
b=>"1110110000",
X=>mulr_4_228);

mulr_1_229<=a_1;
mulc_2_229 : entity work.gfmul
port map(
a=>a_2,
b=>"1100000101",
X=>mulr_2_229);

mulc_3_229 : entity work.gfmul
port map(
a=>a_3,
b=>"1101000011",
X=>mulr_3_229);

mulc_4_229 : entity work.gfmul
port map(
a=>a_4,
b=>"0110111111",
X=>mulr_4_229);

mulr_1_230<=a_1;
mulc_2_230 : entity work.gfmul
port map(
a=>a_2,
b=>"1000000011",
X=>mulr_2_230);

mulc_3_230 : entity work.gfmul
port map(
a=>a_3,
b=>"0100010111",
X=>mulr_3_230);

mulc_4_230 : entity work.gfmul
port map(
a=>a_4,
b=>"0111100011",
X=>mulr_4_230);

mulr_1_231<=a_1;
mulc_2_231 : entity work.gfmul
port map(
a=>a_2,
b=>"0000001111",
X=>mulr_2_231);

mulc_3_231 : entity work.gfmul
port map(
a=>a_3,
b=>"0001010101",
X=>mulr_3_231);

mulc_4_231 : entity work.gfmul
port map(
a=>a_4,
b=>"1100000011",
X=>mulr_4_231);

mulr_1_232<=a_1;
mulc_2_232 : entity work.gfmul
port map(
a=>a_2,
b=>"0000011110",
X=>mulr_2_232);

mulc_3_232 : entity work.gfmul
port map(
a=>a_3,
b=>"0101010100",
X=>mulr_3_232);

mulc_4_232 : entity work.gfmul
port map(
a=>a_4,
b=>"0000101110",
X=>mulr_4_232);

mulr_1_233<=a_1;
mulc_2_233 : entity work.gfmul
port map(
a=>a_2,
b=>"0000111100",
X=>mulr_2_233);

mulc_3_233 : entity work.gfmul
port map(
a=>a_3,
b=>"0101011001",
X=>mulr_3_233);

mulc_4_233 : entity work.gfmul
port map(
a=>a_4,
b=>"0101110000",
X=>mulr_4_233);

mulr_1_234<=a_1;
mulc_2_234 : entity work.gfmul
port map(
a=>a_2,
b=>"0001111000",
X=>mulr_2_234);

mulc_3_234 : entity work.gfmul
port map(
a=>a_3,
b=>"0101101101",
X=>mulr_3_234);

mulc_4_234 : entity work.gfmul
port map(
a=>a_4,
b=>"1110010010",
X=>mulr_4_234);

mulr_1_235<=a_1;
mulc_2_235 : entity work.gfmul
port map(
a=>a_2,
b=>"0011110000",
X=>mulr_2_235);

mulc_3_235 : entity work.gfmul
port map(
a=>a_3,
b=>"0110111101",
X=>mulr_3_235);

mulc_4_235 : entity work.gfmul
port map(
a=>a_4,
b=>"0010101111",
X=>mulr_4_235);

mulr_1_236<=a_1;
mulc_2_236 : entity work.gfmul
port map(
a=>a_2,
b=>"0111100000",
X=>mulr_2_236);

mulc_3_236 : entity work.gfmul
port map(
a=>a_3,
b=>"1011111101",
X=>mulr_3_236);

mulc_4_236 : entity work.gfmul
port map(
a=>a_4,
b=>"0101110001",
X=>mulr_4_236);

mulr_1_237<=a_1;
mulc_2_237 : entity work.gfmul
port map(
a=>a_2,
b=>"1111000000",
X=>mulr_2_237);

mulc_3_237 : entity work.gfmul
port map(
a=>a_3,
b=>"1111100110",
X=>mulr_3_237);

mulc_4_237 : entity work.gfmul
port map(
a=>a_4,
b=>"1110011010",
X=>mulr_4_237);

mulr_1_238<=a_1;
mulc_2_238 : entity work.gfmul
port map(
a=>a_2,
b=>"1110001001",
X=>mulr_2_238);

mulc_3_238 : entity work.gfmul
port map(
a=>a_3,
b=>"1110000011",
X=>mulr_3_238);

mulc_4_238 : entity work.gfmul
port map(
a=>a_4,
b=>"0011101111",
X=>mulr_4_238);

mulr_1_239<=a_1;
mulc_2_239 : entity work.gfmul
port map(
a=>a_2,
b=>"1100011011",
X=>mulr_2_239);

mulc_3_239 : entity work.gfmul
port map(
a=>a_3,
b=>"1000010111",
X=>mulr_3_239);

mulc_4_239 : entity work.gfmul
port map(
a=>a_4,
b=>"1101110001",
X=>mulr_4_239);

mulr_1_240<=a_1;
mulc_2_240 : entity work.gfmul
port map(
a=>a_2,
b=>"1000111111",
X=>mulr_2_240);

mulc_3_240 : entity work.gfmul
port map(
a=>a_3,
b=>"0001001110",
X=>mulr_3_240);

mulc_4_240 : entity work.gfmul
port map(
a=>a_4,
b=>"1110111110",
X=>mulr_4_240);

mulr_1_241<=a_1;
mulc_2_241 : entity work.gfmul
port map(
a=>a_2,
b=>"0001110111",
X=>mulr_2_241);

mulc_3_241 : entity work.gfmul
port map(
a=>a_3,
b=>"0100111000",
X=>mulr_3_241);

mulc_4_241 : entity work.gfmul
port map(
a=>a_4,
b=>"0111001111",
X=>mulr_4_241);

mulr_1_242<=a_1;
mulc_2_242 : entity work.gfmul
port map(
a=>a_2,
b=>"0011101110",
X=>mulr_2_242);

mulc_3_242 : entity work.gfmul
port map(
a=>a_3,
b=>"0011101001",
X=>mulr_3_242);

mulc_4_242 : entity work.gfmul
port map(
a=>a_4,
b=>"1001100011",
X=>mulr_4_242);

mulr_1_243<=a_1;
mulc_2_243 : entity work.gfmul
port map(
a=>a_2,
b=>"0111011100",
X=>mulr_2_243);

mulc_3_243 : entity work.gfmul
port map(
a=>a_3,
b=>"1110100100",
X=>mulr_3_243);

mulc_4_243 : entity work.gfmul
port map(
a=>a_4,
b=>"1100111100",
X=>mulr_4_243);

mulr_1_244<=a_1;
mulc_2_244 : entity work.gfmul
port map(
a=>a_2,
b=>"1110111000",
X=>mulr_2_244);

mulc_3_244 : entity work.gfmul
port map(
a=>a_3,
b=>"1010001011",
X=>mulr_3_244);

mulc_4_244 : entity work.gfmul
port map(
a=>a_4,
b=>"0111010110",
X=>mulr_4_244);

mulr_1_245<=a_1;
mulc_2_245 : entity work.gfmul
port map(
a=>a_2,
b=>"1101111001",
X=>mulr_2_245);

mulc_3_245 : entity work.gfmul
port map(
a=>a_3,
b=>"1000111110",
X=>mulr_3_245);

mulc_4_245 : entity work.gfmul
port map(
a=>a_4,
b=>"1010101011",
X=>mulr_4_245);

mulr_1_246<=a_1;
mulc_2_246 : entity work.gfmul
port map(
a=>a_2,
b=>"1011111011",
X=>mulr_2_246);

mulc_3_246 : entity work.gfmul
port map(
a=>a_3,
b=>"0011101010",
X=>mulr_3_246);

mulc_4_246 : entity work.gfmul
port map(
a=>a_4,
b=>"0101110101",
X=>mulr_4_246);

mulr_1_247<=a_1;
mulc_2_247 : entity work.gfmul
port map(
a=>a_2,
b=>"0111111111",
X=>mulr_2_247);

mulc_3_247 : entity work.gfmul
port map(
a=>a_3,
b=>"1110101000",
X=>mulr_3_247);

mulc_4_247 : entity work.gfmul
port map(
a=>a_4,
b=>"1110111010",
X=>mulr_4_247);

mulr_1_248<=a_1;
mulc_2_248 : entity work.gfmul
port map(
a=>a_2,
b=>"1111111110",
X=>mulr_2_248);

mulc_3_248 : entity work.gfmul
port map(
a=>a_3,
b=>"1010111011",
X=>mulr_3_248);

mulc_4_248 : entity work.gfmul
port map(
a=>a_4,
b=>"0111101111",
X=>mulr_4_248);

mulr_1_249<=a_1;
mulc_2_249 : entity work.gfmul
port map(
a=>a_2,
b=>"1111110101",
X=>mulr_2_249);

mulc_3_249 : entity work.gfmul
port map(
a=>a_3,
b=>"1011111110",
X=>mulr_3_249);

mulc_4_249 : entity work.gfmul
port map(
a=>a_4,
b=>"1101100011",
X=>mulr_4_249);

mulr_1_250<=a_1;
mulc_2_250 : entity work.gfmul
port map(
a=>a_2,
b=>"1111100011",
X=>mulr_2_250);

mulc_3_250 : entity work.gfmul
port map(
a=>a_3,
b=>"1111101010",
X=>mulr_3_250);

mulc_4_250 : entity work.gfmul
port map(
a=>a_4,
b=>"1100101110",
X=>mulr_4_250);

mulr_1_251<=a_1;
mulc_2_251 : entity work.gfmul
port map(
a=>a_2,
b=>"1111001111",
X=>mulr_2_251);

mulc_3_251 : entity work.gfmul
port map(
a=>a_3,
b=>"1110110011",
X=>mulr_3_251);

mulc_4_251 : entity work.gfmul
port map(
a=>a_4,
b=>"0101000110",
X=>mulr_4_251);

mulr_1_252<=a_1;
mulc_2_252 : entity work.gfmul
port map(
a=>a_2,
b=>"1110010111",
X=>mulr_2_252);

mulc_3_252 : entity work.gfmul
port map(
a=>a_3,
b=>"1011010111",
X=>mulr_3_252);

mulc_4_252 : entity work.gfmul
port map(
a=>a_4,
b=>"1000100010",
X=>mulr_4_252);

mulr_1_253<=a_1;
mulc_2_253 : entity work.gfmul
port map(
a=>a_2,
b=>"1100100111",
X=>mulr_2_253);

mulc_3_253 : entity work.gfmul
port map(
a=>a_3,
b=>"1101001110",
X=>mulr_3_253);

mulc_4_253 : entity work.gfmul
port map(
a=>a_4,
b=>"0100110100",
X=>mulr_4_253);

mulr_1_254<=a_1;
mulc_2_254 : entity work.gfmul
port map(
a=>a_2,
b=>"1001000111",
X=>mulr_2_254);

mulc_3_254 : entity work.gfmul
port map(
a=>a_3,
b=>"0100100011",
X=>mulr_3_254);

mulc_4_254 : entity work.gfmul
port map(
a=>a_4,
b=>"0110110010",
X=>mulr_4_254);

mulr_1_255<=a_1;
mulc_2_255 : entity work.gfmul
port map(
a=>a_2,
b=>"0010000111",
X=>mulr_2_255);

mulc_3_255 : entity work.gfmul
port map(
a=>a_3,
b=>"0010000101",
X=>mulr_3_255);

mulc_4_255 : entity work.gfmul
port map(
a=>a_4,
b=>"0110001011",
X=>mulr_4_255);

mulr_1_256<=a_1;
mulc_2_256 : entity work.gfmul
port map(
a=>a_2,
b=>"0100001110",
X=>mulr_2_256);

mulc_3_256 : entity work.gfmul
port map(
a=>a_3,
b=>"1000010100",
X=>mulr_3_256);

mulc_4_256 : entity work.gfmul
port map(
a=>a_4,
b=>"0001000011",
X=>mulr_4_256);

mulr_1_257<=a_1;
mulc_2_257 : entity work.gfmul
port map(
a=>a_2,
b=>"1000011100",
X=>mulr_2_257);

mulc_3_257 : entity work.gfmul
port map(
a=>a_3,
b=>"0001000010",
X=>mulr_3_257);

mulc_4_257 : entity work.gfmul
port map(
a=>a_4,
b=>"1000011000",
X=>mulr_4_257);

mulr_1_258<=a_1;
mulc_2_258 : entity work.gfmul
port map(
a=>a_2,
b=>"0000110001",
X=>mulr_2_258);

mulc_3_258 : entity work.gfmul
port map(
a=>a_3,
b=>"0100001000",
X=>mulr_3_258);

mulc_4_258 : entity work.gfmul
port map(
a=>a_4,
b=>"0011100100",
X=>mulr_4_258);

mulr_1_259<=a_1;
mulc_2_259 : entity work.gfmul
port map(
a=>a_2,
b=>"0001100010",
X=>mulr_2_259);

mulc_3_259 : entity work.gfmul
port map(
a=>a_3,
b=>"0000101001",
X=>mulr_3_259);

mulc_4_259 : entity work.gfmul
port map(
a=>a_4,
b=>"1100101001",
X=>mulr_4_259);

mulr_1_260<=a_1;
mulc_2_260 : entity work.gfmul
port map(
a=>a_2,
b=>"0011000100",
X=>mulr_2_260);

mulc_3_260 : entity work.gfmul
port map(
a=>a_3,
b=>"0010100100",
X=>mulr_3_260);

mulc_4_260 : entity work.gfmul
port map(
a=>a_4,
b=>"0101111110",
X=>mulr_4_260);

mulr_1_261<=a_1;
mulc_2_261 : entity work.gfmul
port map(
a=>a_2,
b=>"0110001000",
X=>mulr_2_261);

mulc_3_261 : entity work.gfmul
port map(
a=>a_3,
b=>"1010010000",
X=>mulr_3_261);

mulc_4_261 : entity work.gfmul
port map(
a=>a_4,
b=>"1111100010",
X=>mulr_4_261);

mulr_1_262<=a_1;
mulc_2_262 : entity work.gfmul
port map(
a=>a_2,
b=>"1100010000",
X=>mulr_2_262);

mulc_3_262 : entity work.gfmul
port map(
a=>a_3,
b=>"1001010010",
X=>mulr_3_262);

mulc_4_262 : entity work.gfmul
port map(
a=>a_4,
b=>"1100101111",
X=>mulr_4_262);

mulr_1_263<=a_1;
mulc_2_263 : entity work.gfmul
port map(
a=>a_2,
b=>"1000101001",
X=>mulr_2_263);

mulc_3_263 : entity work.gfmul
port map(
a=>a_3,
b=>"0101011010",
X=>mulr_3_263);

mulc_4_263 : entity work.gfmul
port map(
a=>a_4,
b=>"0101001110",
X=>mulr_4_263);

mulr_1_264<=a_1;
mulc_2_264 : entity work.gfmul
port map(
a=>a_2,
b=>"0001011011",
X=>mulr_2_264);

mulc_3_264 : entity work.gfmul
port map(
a=>a_3,
b=>"0101100001",
X=>mulr_3_264);

mulc_4_264 : entity work.gfmul
port map(
a=>a_4,
b=>"1001100010",
X=>mulr_4_264);

mulr_1_265<=a_1;
mulc_2_265 : entity work.gfmul
port map(
a=>a_2,
b=>"0010110110",
X=>mulr_2_265);

mulc_3_265 : entity work.gfmul
port map(
a=>a_3,
b=>"0110001101",
X=>mulr_3_265);

mulc_4_265 : entity work.gfmul
port map(
a=>a_4,
b=>"1100110100",
X=>mulr_4_265);

mulr_1_266<=a_1;
mulc_2_266 : entity work.gfmul
port map(
a=>a_2,
b=>"0101101100",
X=>mulr_2_266);

mulc_3_266 : entity work.gfmul
port map(
a=>a_3,
b=>"1000111101",
X=>mulr_3_266);

mulc_4_266 : entity work.gfmul
port map(
a=>a_4,
b=>"0110010110",
X=>mulr_4_266);

mulr_1_267<=a_1;
mulc_2_267 : entity work.gfmul
port map(
a=>a_2,
b=>"1011011000",
X=>mulr_2_267);

mulc_3_267 : entity work.gfmul
port map(
a=>a_3,
b=>"0011100110",
X=>mulr_3_267);

mulc_4_267 : entity work.gfmul
port map(
a=>a_4,
b=>"0010101011",
X=>mulr_4_267);

mulr_1_268<=a_1;
mulc_2_268 : entity work.gfmul
port map(
a=>a_2,
b=>"0110111001",
X=>mulr_2_268);

mulc_3_268 : entity work.gfmul
port map(
a=>a_3,
b=>"1110011000",
X=>mulr_3_268);

mulc_4_268 : entity work.gfmul
port map(
a=>a_4,
b=>"0101010001",
X=>mulr_4_268);

mulr_1_269<=a_1;
mulc_2_269 : entity work.gfmul
port map(
a=>a_2,
b=>"1101110010",
X=>mulr_2_269);

mulc_3_269 : entity work.gfmul
port map(
a=>a_3,
b=>"1001111011",
X=>mulr_3_269);

mulc_4_269 : entity work.gfmul
port map(
a=>a_4,
b=>"1010011010",
X=>mulr_4_269);

mulr_1_270<=a_1;
mulc_2_270 : entity work.gfmul
port map(
a=>a_2,
b=>"1011101101",
X=>mulr_2_270);

mulc_3_270 : entity work.gfmul
port map(
a=>a_3,
b=>"0111111110",
X=>mulr_3_270);

mulc_4_270 : entity work.gfmul
port map(
a=>a_4,
b=>"0011111101",
X=>mulr_4_270);

mulr_1_271<=a_1;
mulc_2_271 : entity work.gfmul
port map(
a=>a_2,
b=>"0111010011",
X=>mulr_2_271);

mulc_3_271 : entity work.gfmul
port map(
a=>a_3,
b=>"1111110001",
X=>mulr_3_271);

mulc_4_271 : entity work.gfmul
port map(
a=>a_4,
b=>"1111100001",
X=>mulr_4_271);

mulr_1_272<=a_1;
mulc_2_272 : entity work.gfmul
port map(
a=>a_2,
b=>"1110100110",
X=>mulr_2_272);

mulc_3_272 : entity work.gfmul
port map(
a=>a_3,
b=>"1111011111",
X=>mulr_3_272);

mulc_4_272 : entity work.gfmul
port map(
a=>a_4,
b=>"1100110111",
X=>mulr_4_272);

mulr_1_273<=a_1;
mulc_2_273 : entity work.gfmul
port map(
a=>a_2,
b=>"1101000101",
X=>mulr_2_273);

mulc_3_273 : entity work.gfmul
port map(
a=>a_3,
b=>"1101100111",
X=>mulr_3_273);

mulc_4_273 : entity work.gfmul
port map(
a=>a_4,
b=>"0110001110",
X=>mulr_4_273);

mulr_1_274<=a_1;
mulc_2_274 : entity work.gfmul
port map(
a=>a_2,
b=>"1010000011",
X=>mulr_2_274);

mulc_3_274 : entity work.gfmul
port map(
a=>a_3,
b=>"0110000111",
X=>mulr_3_274);

mulc_4_274 : entity work.gfmul
port map(
a=>a_4,
b=>"0001101011",
X=>mulr_4_274);

mulr_1_275<=a_1;
mulc_2_275 : entity work.gfmul
port map(
a=>a_2,
b=>"0100001111",
X=>mulr_2_275);

mulc_3_275 : entity work.gfmul
port map(
a=>a_3,
b=>"1000010101",
X=>mulr_3_275);

mulc_4_275 : entity work.gfmul
port map(
a=>a_4,
b=>"1101011000",
X=>mulr_4_275);

mulr_1_276<=a_1;
mulc_2_276 : entity work.gfmul
port map(
a=>a_2,
b=>"1000011110",
X=>mulr_2_276);

mulc_3_276 : entity work.gfmul
port map(
a=>a_3,
b=>"0001000110",
X=>mulr_3_276);

mulc_4_276 : entity work.gfmul
port map(
a=>a_4,
b=>"1011110110",
X=>mulr_4_276);

mulr_1_277<=a_1;
mulc_2_277 : entity work.gfmul
port map(
a=>a_2,
b=>"0000110101",
X=>mulr_2_277);

mulc_3_277 : entity work.gfmul
port map(
a=>a_3,
b=>"0100011000",
X=>mulr_3_277);

mulc_4_277 : entity work.gfmul
port map(
a=>a_4,
b=>"1110011101",
X=>mulr_4_277);

mulr_1_278<=a_1;
mulc_2_278 : entity work.gfmul
port map(
a=>a_2,
b=>"0001101010",
X=>mulr_2_278);

mulc_3_278 : entity work.gfmul
port map(
a=>a_3,
b=>"0001101001",
X=>mulr_3_278);

mulc_4_278 : entity work.gfmul
port map(
a=>a_4,
b=>"0011010111",
X=>mulr_4_278);

mulr_1_279<=a_1;
mulc_2_279 : entity work.gfmul
port map(
a=>a_2,
b=>"0011010100",
X=>mulr_2_279);

mulc_3_279 : entity work.gfmul
port map(
a=>a_3,
b=>"0110100100",
X=>mulr_3_279);

mulc_4_279 : entity work.gfmul
port map(
a=>a_4,
b=>"1010110001",
X=>mulr_4_279);

mulr_1_280<=a_1;
mulc_2_280 : entity work.gfmul
port map(
a=>a_2,
b=>"0110101000",
X=>mulr_2_280);

mulc_3_280 : entity work.gfmul
port map(
a=>a_3,
b=>"1010011001",
X=>mulr_3_280);

mulc_4_280 : entity work.gfmul
port map(
a=>a_4,
b=>"0110100101",
X=>mulr_4_280);

mulr_1_281<=a_1;
mulc_2_281 : entity work.gfmul
port map(
a=>a_2,
b=>"1101010000",
X=>mulr_2_281);

mulc_3_281 : entity work.gfmul
port map(
a=>a_3,
b=>"1001110110",
X=>mulr_3_281);

mulc_4_281 : entity work.gfmul
port map(
a=>a_4,
b=>"0100110011",
X=>mulr_4_281);

mulr_1_282<=a_1;
mulc_2_282 : entity work.gfmul
port map(
a=>a_2,
b=>"1010101001",
X=>mulr_2_282);

mulc_3_282 : entity work.gfmul
port map(
a=>a_3,
b=>"0111001010",
X=>mulr_3_282);

mulc_4_282 : entity work.gfmul
port map(
a=>a_4,
b=>"0110001010",
X=>mulr_4_282);

mulr_1_283<=a_1;
mulc_2_283 : entity work.gfmul
port map(
a=>a_2,
b=>"0101011011",
X=>mulr_2_283);

mulc_3_283 : entity work.gfmul
port map(
a=>a_3,
b=>"1100100001",
X=>mulr_3_283);

mulc_4_283 : entity work.gfmul
port map(
a=>a_4,
b=>"0001001011",
X=>mulr_4_283);

mulr_1_284<=a_1;
mulc_2_284 : entity work.gfmul
port map(
a=>a_2,
b=>"1010110110",
X=>mulr_2_284);

mulc_3_284 : entity work.gfmul
port map(
a=>a_3,
b=>"0010011111",
X=>mulr_3_284);

mulc_4_284 : entity work.gfmul
port map(
a=>a_4,
b=>"1001011000",
X=>mulr_4_284);

mulr_1_285<=a_1;
mulc_2_285 : entity work.gfmul
port map(
a=>a_2,
b=>"0101100101",
X=>mulr_2_285);

mulc_3_285 : entity work.gfmul
port map(
a=>a_3,
b=>"1001111100",
X=>mulr_3_285);

mulc_4_285 : entity work.gfmul
port map(
a=>a_4,
b=>"1011100100",
X=>mulr_4_285);

mulr_1_286<=a_1;
mulc_2_286 : entity work.gfmul
port map(
a=>a_2,
b=>"1011001010",
X=>mulr_2_286);

mulc_3_286 : entity work.gfmul
port map(
a=>a_3,
b=>"0111100010",
X=>mulr_3_286);

mulc_4_286 : entity work.gfmul
port map(
a=>a_4,
b=>"1100001101",
X=>mulr_4_286);

mulr_1_287<=a_1;
mulc_2_287 : entity work.gfmul
port map(
a=>a_2,
b=>"0110011101",
X=>mulr_2_287);

mulc_3_287 : entity work.gfmul
port map(
a=>a_3,
b=>"1110000001",
X=>mulr_3_287);

mulc_4_287 : entity work.gfmul
port map(
a=>a_4,
b=>"0001011110",
X=>mulr_4_287);

mulr_1_288<=a_1;
mulc_2_288 : entity work.gfmul
port map(
a=>a_2,
b=>"1100111010",
X=>mulr_2_288);

mulc_3_288 : entity work.gfmul
port map(
a=>a_3,
b=>"1000011111",
X=>mulr_3_288);

mulc_4_288 : entity work.gfmul
port map(
a=>a_4,
b=>"1011110000",
X=>mulr_4_288);

mulr_1_289<=a_1;
mulc_2_289 : entity work.gfmul
port map(
a=>a_2,
b=>"1001111101",
X=>mulr_2_289);

mulc_3_289 : entity work.gfmul
port map(
a=>a_3,
b=>"0001101110",
X=>mulr_3_289);

mulc_4_289 : entity work.gfmul
port map(
a=>a_4,
b=>"1110101101",
X=>mulr_4_289);

mulr_1_290<=a_1;
mulc_2_290 : entity work.gfmul
port map(
a=>a_2,
b=>"0011110011",
X=>mulr_2_290);

mulc_3_290 : entity work.gfmul
port map(
a=>a_3,
b=>"0110111000",
X=>mulr_3_290);

mulc_4_290 : entity work.gfmul
port map(
a=>a_4,
b=>"0101010111",
X=>mulr_4_290);

mulr_1_291<=a_1;
mulc_2_291 : entity work.gfmul
port map(
a=>a_2,
b=>"0111100110",
X=>mulr_2_291);

mulc_3_291 : entity work.gfmul
port map(
a=>a_3,
b=>"1011101001",
X=>mulr_3_291);

mulc_4_291 : entity work.gfmul
port map(
a=>a_4,
b=>"1010101010",
X=>mulr_4_291);

mulr_1_292<=a_1;
mulc_2_292 : entity work.gfmul
port map(
a=>a_2,
b=>"1111001100",
X=>mulr_2_292);

mulc_3_292 : entity work.gfmul
port map(
a=>a_3,
b=>"1110110110",
X=>mulr_3_292);

mulc_4_292 : entity work.gfmul
port map(
a=>a_4,
b=>"0101111101",
X=>mulr_4_292);

mulr_1_293<=a_1;
mulc_2_293 : entity work.gfmul
port map(
a=>a_2,
b=>"1110010001",
X=>mulr_2_293);

mulc_3_293 : entity work.gfmul
port map(
a=>a_3,
b=>"1011000011",
X=>mulr_3_293);

mulc_4_293 : entity work.gfmul
port map(
a=>a_4,
b=>"1111111010",
X=>mulr_4_293);

mulr_1_294<=a_1;
mulc_2_294 : entity work.gfmul
port map(
a=>a_2,
b=>"1100101011",
X=>mulr_2_294);

mulc_3_294 : entity work.gfmul
port map(
a=>a_3,
b=>"1100011110",
X=>mulr_3_294);

mulc_4_294 : entity work.gfmul
port map(
a=>a_4,
b=>"1111101111",
X=>mulr_4_294);

mulr_1_295<=a_1;
mulc_2_295 : entity work.gfmul
port map(
a=>a_2,
b=>"1001011111",
X=>mulr_2_295);

mulc_3_295 : entity work.gfmul
port map(
a=>a_3,
b=>"0001100011",
X=>mulr_3_295);

mulc_4_295 : entity work.gfmul
port map(
a=>a_4,
b=>"1101000111",
X=>mulr_4_295);

mulr_1_296<=a_1;
mulc_2_296 : entity work.gfmul
port map(
a=>a_2,
b=>"0010110111",
X=>mulr_2_296);

mulc_3_296 : entity work.gfmul
port map(
a=>a_3,
b=>"0110001100",
X=>mulr_3_296);

mulc_4_296 : entity work.gfmul
port map(
a=>a_4,
b=>"1000001110",
X=>mulr_4_296);

mulr_1_297<=a_1;
mulc_2_297 : entity work.gfmul
port map(
a=>a_2,
b=>"0101101110",
X=>mulr_2_297);

mulc_3_297 : entity work.gfmul
port map(
a=>a_3,
b=>"1000111001",
X=>mulr_3_297);

mulc_4_297 : entity work.gfmul
port map(
a=>a_4,
b=>"0001010100",
X=>mulr_4_297);

mulr_1_298<=a_1;
mulc_2_298 : entity work.gfmul
port map(
a=>a_2,
b=>"1011011100",
X=>mulr_2_298);

mulc_3_298 : entity work.gfmul
port map(
a=>a_3,
b=>"0011110110",
X=>mulr_3_298);

mulc_4_298 : entity work.gfmul
port map(
a=>a_4,
b=>"1010100000",
X=>mulr_4_298);

mulr_1_299<=a_1;
mulc_2_299 : entity work.gfmul
port map(
a=>a_2,
b=>"0110110001",
X=>mulr_2_299);

mulc_3_299 : entity work.gfmul
port map(
a=>a_3,
b=>"1111011000",
X=>mulr_3_299);

mulc_4_299 : entity work.gfmul
port map(
a=>a_4,
b=>"0100101101",
X=>mulr_4_299);

mulr_1_300<=a_1;
mulc_2_300 : entity work.gfmul
port map(
a=>a_2,
b=>"1101100010",
X=>mulr_2_300);

mulc_3_300 : entity work.gfmul
port map(
a=>a_3,
b=>"1101111011",
X=>mulr_3_300);

mulc_4_300 : entity work.gfmul
port map(
a=>a_4,
b=>"0101111010",
X=>mulr_4_300);

mulr_1_301<=a_1;
mulc_2_301 : entity work.gfmul
port map(
a=>a_2,
b=>"1011001101",
X=>mulr_2_301);

mulc_3_301 : entity work.gfmul
port map(
a=>a_3,
b=>"0111110111",
X=>mulr_3_301);

mulc_4_301 : entity work.gfmul
port map(
a=>a_4,
b=>"1111000010",
X=>mulr_4_301);

mulr_1_302<=a_1;
mulc_2_302 : entity work.gfmul
port map(
a=>a_2,
b=>"0110010011",
X=>mulr_2_302);

mulc_3_302 : entity work.gfmul
port map(
a=>a_3,
b=>"1111010101",
X=>mulr_3_302);

mulc_4_302 : entity work.gfmul
port map(
a=>a_4,
b=>"1000101111",
X=>mulr_4_302);

mulr_1_303<=a_1;
mulc_2_303 : entity work.gfmul
port map(
a=>a_2,
b=>"1100100110",
X=>mulr_2_303);

mulc_3_303 : entity work.gfmul
port map(
a=>a_3,
b=>"1101001111",
X=>mulr_3_303);

mulc_4_303 : entity work.gfmul
port map(
a=>a_4,
b=>"0101011100",
X=>mulr_4_303);

mulr_1_304<=a_1;
mulc_2_304 : entity work.gfmul
port map(
a=>a_2,
b=>"1001000101",
X=>mulr_2_304);

mulc_3_304 : entity work.gfmul
port map(
a=>a_3,
b=>"0100100111",
X=>mulr_3_304);

mulc_4_304 : entity work.gfmul
port map(
a=>a_4,
b=>"1011110010",
X=>mulr_4_304);

mulr_1_305<=a_1;
mulc_2_305 : entity work.gfmul
port map(
a=>a_2,
b=>"0010000011",
X=>mulr_2_305);

mulc_3_305 : entity work.gfmul
port map(
a=>a_3,
b=>"0010010101",
X=>mulr_3_305);

mulc_4_305 : entity work.gfmul
port map(
a=>a_4,
b=>"1110111101",
X=>mulr_4_305);

mulr_1_306<=a_1;
mulc_2_306 : entity work.gfmul
port map(
a=>a_2,
b=>"0100000110",
X=>mulr_2_306);

mulc_3_306 : entity work.gfmul
port map(
a=>a_3,
b=>"1001010100",
X=>mulr_3_306);

mulc_4_306 : entity work.gfmul
port map(
a=>a_4,
b=>"0111010111",
X=>mulr_4_306);

mulr_1_307<=a_1;
mulc_2_307 : entity work.gfmul
port map(
a=>a_2,
b=>"1000001100",
X=>mulr_2_307);

mulc_3_307 : entity work.gfmul
port map(
a=>a_3,
b=>"0101000010",
X=>mulr_3_307);

mulc_4_307 : entity work.gfmul
port map(
a=>a_4,
b=>"1010100011",
X=>mulr_4_307);

mulr_1_308<=a_1;
mulc_2_308 : entity work.gfmul
port map(
a=>a_2,
b=>"0000010001",
X=>mulr_2_308);

mulc_3_308 : entity work.gfmul
port map(
a=>a_3,
b=>"0100000001",
X=>mulr_3_308);

mulc_4_308 : entity work.gfmul
port map(
a=>a_4,
b=>"0100110101",
X=>mulr_4_308);

mulr_1_309<=a_1;
mulc_2_309 : entity work.gfmul
port map(
a=>a_2,
b=>"0000100010",
X=>mulr_2_309);

mulc_3_309 : entity work.gfmul
port map(
a=>a_3,
b=>"0000001101",
X=>mulr_3_309);

mulc_4_309 : entity work.gfmul
port map(
a=>a_4,
b=>"0110111010",
X=>mulr_4_309);

mulr_1_310<=a_1;
mulc_2_310 : entity work.gfmul
port map(
a=>a_2,
b=>"0001000100",
X=>mulr_2_310);

mulc_3_310 : entity work.gfmul
port map(
a=>a_3,
b=>"0000110100",
X=>mulr_3_310);

mulc_4_310 : entity work.gfmul
port map(
a=>a_4,
b=>"0111001011",
X=>mulr_4_310);

mulr_1_311<=a_1;
mulc_2_311 : entity work.gfmul
port map(
a=>a_2,
b=>"0010001000",
X=>mulr_2_311);

mulc_3_311 : entity work.gfmul
port map(
a=>a_3,
b=>"0011010000",
X=>mulr_3_311);

mulc_4_311 : entity work.gfmul
port map(
a=>a_4,
b=>"1001000011",
X=>mulr_4_311);

mulr_1_312<=a_1;
mulc_2_312 : entity work.gfmul
port map(
a=>a_2,
b=>"0100010000",
X=>mulr_2_312);

mulc_3_312 : entity work.gfmul
port map(
a=>a_3,
b=>"1101000000",
X=>mulr_3_312);

mulc_4_312 : entity work.gfmul
port map(
a=>a_4,
b=>"1000111100",
X=>mulr_4_312);

mulr_1_313<=a_1;
mulc_2_313 : entity work.gfmul
port map(
a=>a_2,
b=>"1000100000",
X=>mulr_2_313);

mulc_3_313 : entity work.gfmul
port map(
a=>a_3,
b=>"0100011011",
X=>mulr_3_313);

mulc_4_313 : entity work.gfmul
port map(
a=>a_4,
b=>"0111000100",
X=>mulr_4_313);

mulr_1_314<=a_1;
mulc_2_314 : entity work.gfmul
port map(
a=>a_2,
b=>"0001001001",
X=>mulr_2_314);

mulc_3_314 : entity work.gfmul
port map(
a=>a_3,
b=>"0001100101",
X=>mulr_3_314);

mulc_4_314 : entity work.gfmul
port map(
a=>a_4,
b=>"1000111011",
X=>mulr_4_314);

mulr_1_315<=a_1;
mulc_2_315 : entity work.gfmul
port map(
a=>a_2,
b=>"0010010010",
X=>mulr_2_315);

mulc_3_315 : entity work.gfmul
port map(
a=>a_3,
b=>"0110010100",
X=>mulr_3_315);

mulc_4_315 : entity work.gfmul
port map(
a=>a_4,
b=>"0111111100",
X=>mulr_4_315);

mulr_1_316<=a_1;
mulc_2_316 : entity work.gfmul
port map(
a=>a_2,
b=>"0100100100",
X=>mulr_2_316);

mulc_3_316 : entity work.gfmul
port map(
a=>a_3,
b=>"1001011001",
X=>mulr_3_316);

mulc_4_316 : entity work.gfmul
port map(
a=>a_4,
b=>"1111111011",
X=>mulr_4_316);

mulr_1_317<=a_1;
mulc_2_317 : entity work.gfmul
port map(
a=>a_2,
b=>"1001001000",
X=>mulr_2_317);

mulc_3_317 : entity work.gfmul
port map(
a=>a_3,
b=>"0101110110",
X=>mulr_3_317);

mulc_4_317 : entity work.gfmul
port map(
a=>a_4,
b=>"1111100111",
X=>mulr_4_317);

mulr_1_318<=a_1;
mulc_2_318 : entity work.gfmul
port map(
a=>a_2,
b=>"0010011001",
X=>mulr_2_318);

mulc_3_318 : entity work.gfmul
port map(
a=>a_3,
b=>"0111010001",
X=>mulr_3_318);

mulc_4_318 : entity work.gfmul
port map(
a=>a_4,
b=>"1100000111",
X=>mulr_4_318);

mulr_1_319<=a_1;
mulc_2_319 : entity work.gfmul
port map(
a=>a_2,
b=>"0100110010",
X=>mulr_2_319);

mulc_3_319 : entity work.gfmul
port map(
a=>a_3,
b=>"1101001101",
X=>mulr_3_319);

mulc_4_319 : entity work.gfmul
port map(
a=>a_4,
b=>"0000001110",
X=>mulr_4_319);

mulr_1_320<=a_1;
mulc_2_320 : entity work.gfmul
port map(
a=>a_2,
b=>"1001100100",
X=>mulr_2_320);

mulc_3_320 : entity work.gfmul
port map(
a=>a_3,
b=>"0100101111",
X=>mulr_3_320);

mulc_4_320 : entity work.gfmul
port map(
a=>a_4,
b=>"0001110000",
X=>mulr_4_320);

mulr_1_321<=a_1;
mulc_2_321 : entity work.gfmul
port map(
a=>a_2,
b=>"0011000001",
X=>mulr_2_321);

mulc_3_321 : entity work.gfmul
port map(
a=>a_3,
b=>"0010110101",
X=>mulr_3_321);

mulc_4_321 : entity work.gfmul
port map(
a=>a_4,
b=>"1110000000",
X=>mulr_4_321);

mulr_1_322<=a_1;
mulc_2_322 : entity work.gfmul
port map(
a=>a_2,
b=>"0110000010",
X=>mulr_2_322);

mulc_3_322 : entity work.gfmul
port map(
a=>a_3,
b=>"1011010100",
X=>mulr_3_322);

mulc_4_322 : entity work.gfmul
port map(
a=>a_4,
b=>"0000111111",
X=>mulr_4_322);

mulr_1_323<=a_1;
mulc_2_323 : entity work.gfmul
port map(
a=>a_2,
b=>"1100000100",
X=>mulr_2_323);

mulc_3_323 : entity work.gfmul
port map(
a=>a_3,
b=>"1101000010",
X=>mulr_3_323);

mulc_4_323 : entity work.gfmul
port map(
a=>a_4,
b=>"0111111000",
X=>mulr_4_323);

mulr_1_324<=a_1;
mulc_2_324 : entity work.gfmul
port map(
a=>a_2,
b=>"1000000001",
X=>mulr_2_324);

mulc_3_324 : entity work.gfmul
port map(
a=>a_3,
b=>"0100010011",
X=>mulr_3_324);

mulc_4_324 : entity work.gfmul
port map(
a=>a_4,
b=>"1111011011",
X=>mulr_4_324);

mulr_1_325<=a_1;
mulc_2_325 : entity work.gfmul
port map(
a=>a_2,
b=>"0000001011",
X=>mulr_2_325);

mulc_3_325 : entity work.gfmul
port map(
a=>a_3,
b=>"0001000101",
X=>mulr_3_325);

mulc_4_325 : entity work.gfmul
port map(
a=>a_4,
b=>"1011100111",
X=>mulr_4_325);

mulr_1_326<=a_1;
mulc_2_326 : entity work.gfmul
port map(
a=>a_2,
b=>"0000010110",
X=>mulr_2_326);

mulc_3_326 : entity work.gfmul
port map(
a=>a_3,
b=>"0100010100",
X=>mulr_3_326);

mulc_4_326 : entity work.gfmul
port map(
a=>a_4,
b=>"1100010101",
X=>mulr_4_326);

mulr_1_327<=a_1;
mulc_2_327 : entity work.gfmul
port map(
a=>a_2,
b=>"0000101100",
X=>mulr_2_327);

mulc_3_327 : entity work.gfmul
port map(
a=>a_3,
b=>"0001011001",
X=>mulr_3_327);

mulc_4_327 : entity work.gfmul
port map(
a=>a_4,
b=>"0010011110",
X=>mulr_4_327);

mulr_1_328<=a_1;
mulc_2_328 : entity work.gfmul
port map(
a=>a_2,
b=>"0001011000",
X=>mulr_2_328);

mulc_3_328 : entity work.gfmul
port map(
a=>a_3,
b=>"0101100100",
X=>mulr_3_328);

mulc_4_328 : entity work.gfmul
port map(
a=>a_4,
b=>"0011111001",
X=>mulr_4_328);

mulr_1_329<=a_1;
mulc_2_329 : entity work.gfmul
port map(
a=>a_2,
b=>"0010110000",
X=>mulr_2_329);

mulc_3_329 : entity work.gfmul
port map(
a=>a_3,
b=>"0110011001",
X=>mulr_3_329);

mulc_4_329 : entity work.gfmul
port map(
a=>a_4,
b=>"1111000001",
X=>mulr_4_329);

mulr_1_330<=a_1;
mulc_2_330 : entity work.gfmul
port map(
a=>a_2,
b=>"0101100000",
X=>mulr_2_330);

mulc_3_330 : entity work.gfmul
port map(
a=>a_3,
b=>"1001101101",
X=>mulr_3_330);

mulc_4_330 : entity work.gfmul
port map(
a=>a_4,
b=>"1000110111",
X=>mulr_4_330);

mulr_1_331<=a_1;
mulc_2_331 : entity work.gfmul
port map(
a=>a_2,
b=>"1011000000",
X=>mulr_2_331);

mulc_3_331 : entity work.gfmul
port map(
a=>a_3,
b=>"0110100110",
X=>mulr_3_331);

mulc_4_331 : entity work.gfmul
port map(
a=>a_4,
b=>"0110011100",
X=>mulr_4_331);

mulr_1_332<=a_1;
mulc_2_332 : entity work.gfmul
port map(
a=>a_2,
b=>"0110001001",
X=>mulr_2_332);

mulc_3_332 : entity work.gfmul
port map(
a=>a_3,
b=>"1010010001",
X=>mulr_3_332);

mulc_4_332 : entity work.gfmul
port map(
a=>a_4,
b=>"0011111011",
X=>mulr_4_332);

mulr_1_333<=a_1;
mulc_2_333 : entity work.gfmul
port map(
a=>a_2,
b=>"1100010010",
X=>mulr_2_333);

mulc_3_333 : entity work.gfmul
port map(
a=>a_3,
b=>"1001010110",
X=>mulr_3_333);

mulc_4_333 : entity work.gfmul
port map(
a=>a_4,
b=>"1111010001",
X=>mulr_4_333);

mulr_1_334<=a_1;
mulc_2_334 : entity work.gfmul
port map(
a=>a_2,
b=>"1000101101",
X=>mulr_2_334);

mulc_3_334 : entity work.gfmul
port map(
a=>a_3,
b=>"0101001010",
X=>mulr_3_334);

mulc_4_334 : entity work.gfmul
port map(
a=>a_4,
b=>"1010110111",
X=>mulr_4_334);

mulr_1_335<=a_1;
mulc_2_335 : entity work.gfmul
port map(
a=>a_2,
b=>"0001010011",
X=>mulr_2_335);

mulc_3_335 : entity work.gfmul
port map(
a=>a_3,
b=>"0100100001",
X=>mulr_3_335);

mulc_4_335 : entity work.gfmul
port map(
a=>a_4,
b=>"0110010101",
X=>mulr_4_335);

mulr_1_336<=a_1;
mulc_2_336 : entity work.gfmul
port map(
a=>a_2,
b=>"0010100110",
X=>mulr_2_336);

mulc_3_336 : entity work.gfmul
port map(
a=>a_3,
b=>"0010001101",
X=>mulr_3_336);

mulc_4_336 : entity work.gfmul
port map(
a=>a_4,
b=>"0010110011",
X=>mulr_4_336);

mulr_1_337<=a_1;
mulc_2_337 : entity work.gfmul
port map(
a=>a_2,
b=>"0101001100",
X=>mulr_2_337);

mulc_3_337 : entity work.gfmul
port map(
a=>a_3,
b=>"1000110100",
X=>mulr_3_337);

mulc_4_337 : entity work.gfmul
port map(
a=>a_4,
b=>"0110010001",
X=>mulr_4_337);

mulr_1_338<=a_1;
mulc_2_338 : entity work.gfmul
port map(
a=>a_2,
b=>"1010011000",
X=>mulr_2_338);

mulc_3_338 : entity work.gfmul
port map(
a=>a_3,
b=>"0011000010",
X=>mulr_3_338);

mulc_4_338 : entity work.gfmul
port map(
a=>a_4,
b=>"0010010011",
X=>mulr_4_338);

mulr_1_339<=a_1;
mulc_2_339 : entity work.gfmul
port map(
a=>a_2,
b=>"0100111001",
X=>mulr_2_339);

mulc_3_339 : entity work.gfmul
port map(
a=>a_3,
b=>"1100001000",
X=>mulr_3_339);

mulc_4_339 : entity work.gfmul
port map(
a=>a_4,
b=>"0010010001",
X=>mulr_4_339);

mulr_1_340<=a_1;
mulc_2_340 : entity work.gfmul
port map(
a=>a_2,
b=>"1001110010",
X=>mulr_2_340);

mulc_3_340 : entity work.gfmul
port map(
a=>a_3,
b=>"0000111011",
X=>mulr_3_340);

mulc_4_340 : entity work.gfmul
port map(
a=>a_4,
b=>"0010000001",
X=>mulr_4_340);

mulr_1_341<=a_1;
mulc_2_341 : entity work.gfmul
port map(
a=>a_2,
b=>"0011101101",
X=>mulr_2_341);

mulc_3_341 : entity work.gfmul
port map(
a=>a_3,
b=>"0011101100",
X=>mulr_3_341);

mulc_4_341 : entity work.gfmul
port map(
a=>a_4,
b=>"0000000001",
X=>mulr_4_341);

mulr_1_342<=a_1;
mulc_2_342 : entity work.gfmul
port map(
a=>a_2,
b=>"0111011010",
X=>mulr_2_342);

mulc_3_342 : entity work.gfmul
port map(
a=>a_3,
b=>"1110110000",
X=>mulr_3_342);

mulc_4_342 : entity work.gfmul
port map(
a=>a_4,
b=>"0000001000",
X=>mulr_4_342);

mulr_1_343<=a_1;
mulc_2_343 : entity work.gfmul
port map(
a=>a_2,
b=>"1110110100",
X=>mulr_2_343);

mulc_3_343 : entity work.gfmul
port map(
a=>a_3,
b=>"1011011011",
X=>mulr_3_343);

mulc_4_343 : entity work.gfmul
port map(
a=>a_4,
b=>"0001000000",
X=>mulr_4_343);

mulr_1_344<=a_1;
mulc_2_344 : entity work.gfmul
port map(
a=>a_2,
b=>"1101100001",
X=>mulr_2_344);

mulc_3_344 : entity work.gfmul
port map(
a=>a_3,
b=>"1101111110",
X=>mulr_3_344);

mulc_4_344 : entity work.gfmul
port map(
a=>a_4,
b=>"1000000000",
X=>mulr_4_344);

mulr_1_345<=a_1;
mulc_2_345 : entity work.gfmul
port map(
a=>a_2,
b=>"1011001011",
X=>mulr_2_345);

mulc_3_345 : entity work.gfmul
port map(
a=>a_3,
b=>"0111100011",
X=>mulr_3_345);

mulc_4_345 : entity work.gfmul
port map(
a=>a_4,
b=>"0000100100",
X=>mulr_4_345);

mulr_1_346<=a_1;
mulc_2_346 : entity work.gfmul
port map(
a=>a_2,
b=>"0110011111",
X=>mulr_2_346);

mulc_3_346 : entity work.gfmul
port map(
a=>a_3,
b=>"1110000101",
X=>mulr_3_346);

mulc_4_346 : entity work.gfmul
port map(
a=>a_4,
b=>"0100100000",
X=>mulr_4_346);

mulr_1_347<=a_1;
mulc_2_347 : entity work.gfmul
port map(
a=>a_2,
b=>"1100111110",
X=>mulr_2_347);

mulc_3_347 : entity work.gfmul
port map(
a=>a_3,
b=>"1000001111",
X=>mulr_3_347);

mulc_4_347 : entity work.gfmul
port map(
a=>a_4,
b=>"0100010010",
X=>mulr_4_347);

mulr_1_348<=a_1;
mulc_2_348 : entity work.gfmul
port map(
a=>a_2,
b=>"1001110101",
X=>mulr_2_348);

mulc_3_348 : entity work.gfmul
port map(
a=>a_3,
b=>"0000101110",
X=>mulr_3_348);

mulc_4_348 : entity work.gfmul
port map(
a=>a_4,
b=>"0010000010",
X=>mulr_4_348);

mulr_1_349<=a_1;
mulc_2_349 : entity work.gfmul
port map(
a=>a_2,
b=>"0011100011",
X=>mulr_2_349);

mulc_3_349 : entity work.gfmul
port map(
a=>a_3,
b=>"0010111000",
X=>mulr_3_349);

mulc_4_349 : entity work.gfmul
port map(
a=>a_4,
b=>"0000011001",
X=>mulr_4_349);

mulr_1_350<=a_1;
mulc_2_350 : entity work.gfmul
port map(
a=>a_2,
b=>"0111000110",
X=>mulr_2_350);

mulc_3_350 : entity work.gfmul
port map(
a=>a_3,
b=>"1011100000",
X=>mulr_3_350);

mulc_4_350 : entity work.gfmul
port map(
a=>a_4,
b=>"0011001000",
X=>mulr_4_350);

mulr_1_351<=a_1;
mulc_2_351 : entity work.gfmul
port map(
a=>a_2,
b=>"1110001100",
X=>mulr_2_351);

mulc_3_351 : entity work.gfmul
port map(
a=>a_3,
b=>"1110010010",
X=>mulr_3_351);

mulc_4_351 : entity work.gfmul
port map(
a=>a_4,
b=>"1001001001",
X=>mulr_4_351);

mulr_1_352<=a_1;
mulc_2_352 : entity work.gfmul
port map(
a=>a_2,
b=>"1100010001",
X=>mulr_2_352);

mulc_3_352 : entity work.gfmul
port map(
a=>a_3,
b=>"1001010011",
X=>mulr_3_352);

mulc_4_352 : entity work.gfmul
port map(
a=>a_4,
b=>"1001101100",
X=>mulr_4_352);

mulr_1_353<=a_1;
mulc_2_353 : entity work.gfmul
port map(
a=>a_2,
b=>"1000101011",
X=>mulr_2_353);

mulc_3_353 : entity work.gfmul
port map(
a=>a_3,
b=>"0101011110",
X=>mulr_3_353);

mulc_4_353 : entity work.gfmul
port map(
a=>a_4,
b=>"1101000100",
X=>mulr_4_353);

mulr_1_354<=a_1;
mulc_2_354 : entity work.gfmul
port map(
a=>a_2,
b=>"0001011111",
X=>mulr_2_354);

mulc_3_354 : entity work.gfmul
port map(
a=>a_3,
b=>"0101110001",
X=>mulr_3_354);

mulc_4_354 : entity work.gfmul
port map(
a=>a_4,
b=>"1000010110",
X=>mulr_4_354);

mulr_1_355<=a_1;
mulc_2_355 : entity work.gfmul
port map(
a=>a_2,
b=>"0010111110",
X=>mulr_2_355);

mulc_3_355 : entity work.gfmul
port map(
a=>a_3,
b=>"0111001101",
X=>mulr_3_355);

mulc_4_355 : entity work.gfmul
port map(
a=>a_4,
b=>"0010010100",
X=>mulr_4_355);

mulr_1_356<=a_1;
mulc_2_356 : entity work.gfmul
port map(
a=>a_2,
b=>"0101111100",
X=>mulr_2_356);

mulc_3_356 : entity work.gfmul
port map(
a=>a_3,
b=>"1100111101",
X=>mulr_3_356);

mulc_4_356 : entity work.gfmul
port map(
a=>a_4,
b=>"0010101001",
X=>mulr_4_356);

mulr_1_357<=a_1;
mulc_2_357 : entity work.gfmul
port map(
a=>a_2,
b=>"1011111000",
X=>mulr_2_357);

mulc_3_357 : entity work.gfmul
port map(
a=>a_3,
b=>"0011101111",
X=>mulr_3_357);

mulc_4_357 : entity work.gfmul
port map(
a=>a_4,
b=>"0101000001",
X=>mulr_4_357);

mulr_1_358<=a_1;
mulc_2_358 : entity work.gfmul
port map(
a=>a_2,
b=>"0111111001",
X=>mulr_2_358);

mulc_3_358 : entity work.gfmul
port map(
a=>a_3,
b=>"1110111100",
X=>mulr_3_358);

mulc_4_358 : entity work.gfmul
port map(
a=>a_4,
b=>"1000011010",
X=>mulr_4_358);

mulr_1_359<=a_1;
mulc_2_359 : entity work.gfmul
port map(
a=>a_2,
b=>"1111110010",
X=>mulr_2_359);

mulc_3_359 : entity work.gfmul
port map(
a=>a_3,
b=>"1011101011",
X=>mulr_3_359);

mulc_4_359 : entity work.gfmul
port map(
a=>a_4,
b=>"0011110100",
X=>mulr_4_359);

mulr_1_360<=a_1;
mulc_2_360 : entity work.gfmul
port map(
a=>a_2,
b=>"1111101101",
X=>mulr_2_360);

mulc_3_360 : entity work.gfmul
port map(
a=>a_3,
b=>"1110111110",
X=>mulr_3_360);

mulc_4_360 : entity work.gfmul
port map(
a=>a_4,
b=>"1110101001",
X=>mulr_4_360);

mulr_1_361<=a_1;
mulc_2_361 : entity work.gfmul
port map(
a=>a_2,
b=>"1111010011",
X=>mulr_2_361);

mulc_3_361 : entity work.gfmul
port map(
a=>a_3,
b=>"1011100011",
X=>mulr_3_361);

mulc_4_361 : entity work.gfmul
port map(
a=>a_4,
b=>"0101110111",
X=>mulr_4_361);

mulr_1_362<=a_1;
mulc_2_362 : entity work.gfmul
port map(
a=>a_2,
b=>"1110101111",
X=>mulr_2_362);

mulc_3_362 : entity work.gfmul
port map(
a=>a_3,
b=>"1110011110",
X=>mulr_3_362);

mulc_4_362 : entity work.gfmul
port map(
a=>a_4,
b=>"1110101010",
X=>mulr_4_362);

mulr_1_363<=a_1;
mulc_2_363 : entity work.gfmul
port map(
a=>a_2,
b=>"1101010111",
X=>mulr_2_363);

mulc_3_363 : entity work.gfmul
port map(
a=>a_3,
b=>"1001100011",
X=>mulr_3_363);

mulc_4_363 : entity work.gfmul
port map(
a=>a_4,
b=>"0101101111",
X=>mulr_4_363);

mulr_1_364<=a_1;
mulc_2_364 : entity work.gfmul
port map(
a=>a_2,
b=>"1010100111",
X=>mulr_2_364);

mulc_3_364 : entity work.gfmul
port map(
a=>a_3,
b=>"0110011110",
X=>mulr_3_364);

mulc_4_364 : entity work.gfmul
port map(
a=>a_4,
b=>"1101101010",
X=>mulr_4_364);

mulr_1_365<=a_1;
mulc_2_365 : entity work.gfmul
port map(
a=>a_2,
b=>"0101000111",
X=>mulr_2_365);

mulc_3_365 : entity work.gfmul
port map(
a=>a_3,
b=>"1001110001",
X=>mulr_3_365);

mulc_4_365 : entity work.gfmul
port map(
a=>a_4,
b=>"1101100110",
X=>mulr_4_365);

mulr_1_366<=a_1;
mulc_2_366 : entity work.gfmul
port map(
a=>a_2,
b=>"1010001110",
X=>mulr_2_366);

mulc_3_366 : entity work.gfmul
port map(
a=>a_3,
b=>"0111010110",
X=>mulr_3_366);

mulc_4_366 : entity work.gfmul
port map(
a=>a_4,
b=>"1100000110",
X=>mulr_4_366);

mulr_1_367<=a_1;
mulc_2_367 : entity work.gfmul
port map(
a=>a_2,
b=>"0100010101",
X=>mulr_2_367);

mulc_3_367 : entity work.gfmul
port map(
a=>a_3,
b=>"1101010001",
X=>mulr_3_367);

mulc_4_367 : entity work.gfmul
port map(
a=>a_4,
b=>"0000000110",
X=>mulr_4_367);

mulr_1_368<=a_1;
mulc_2_368 : entity work.gfmul
port map(
a=>a_2,
b=>"1000101010",
X=>mulr_2_368);

mulc_3_368 : entity work.gfmul
port map(
a=>a_3,
b=>"0101011111",
X=>mulr_3_368);

mulc_4_368 : entity work.gfmul
port map(
a=>a_4,
b=>"0000110000",
X=>mulr_4_368);

mulr_1_369<=a_1;
mulc_2_369 : entity work.gfmul
port map(
a=>a_2,
b=>"0001011101",
X=>mulr_2_369);

mulc_3_369 : entity work.gfmul
port map(
a=>a_3,
b=>"0101110101",
X=>mulr_3_369);

mulc_4_369 : entity work.gfmul
port map(
a=>a_4,
b=>"0110000000",
X=>mulr_4_369);

mulr_1_370<=a_1;
mulc_2_370 : entity work.gfmul
port map(
a=>a_2,
b=>"0010111010",
X=>mulr_2_370);

mulc_3_370 : entity work.gfmul
port map(
a=>a_3,
b=>"0111011101",
X=>mulr_3_370);

mulc_4_370 : entity work.gfmul
port map(
a=>a_4,
b=>"0000011011",
X=>mulr_4_370);

mulr_1_371<=a_1;
mulc_2_371 : entity work.gfmul
port map(
a=>a_2,
b=>"0101110100",
X=>mulr_2_371);

mulc_3_371 : entity work.gfmul
port map(
a=>a_3,
b=>"1101111101",
X=>mulr_3_371);

mulc_4_371 : entity work.gfmul
port map(
a=>a_4,
b=>"0011011000",
X=>mulr_4_371);

mulr_1_372<=a_1;
mulc_2_372 : entity work.gfmul
port map(
a=>a_2,
b=>"1011101000",
X=>mulr_2_372);

mulc_3_372 : entity work.gfmul
port map(
a=>a_3,
b=>"0111101111",
X=>mulr_3_372);

mulc_4_372 : entity work.gfmul
port map(
a=>a_4,
b=>"1011001001",
X=>mulr_4_372);

mulr_1_373<=a_1;
mulc_2_373 : entity work.gfmul
port map(
a=>a_2,
b=>"0111011001",
X=>mulr_2_373);

mulc_3_373 : entity work.gfmul
port map(
a=>a_3,
b=>"1110110101",
X=>mulr_3_373);

mulc_4_373 : entity work.gfmul
port map(
a=>a_4,
b=>"1001100101",
X=>mulr_4_373);

mulr_1_374<=a_1;
mulc_2_374 : entity work.gfmul
port map(
a=>a_2,
b=>"1110110010",
X=>mulr_2_374);

mulc_3_374 : entity work.gfmul
port map(
a=>a_3,
b=>"1011001111",
X=>mulr_3_374);

mulc_4_374 : entity work.gfmul
port map(
a=>a_4,
b=>"1100001100",
X=>mulr_4_374);

mulr_1_375<=a_1;
mulc_2_375 : entity work.gfmul
port map(
a=>a_2,
b=>"1101101101",
X=>mulr_2_375);

mulc_3_375 : entity work.gfmul
port map(
a=>a_3,
b=>"1100101110",
X=>mulr_3_375);

mulc_4_375 : entity work.gfmul
port map(
a=>a_4,
b=>"0001010110",
X=>mulr_4_375);

mulr_1_376<=a_1;
mulc_2_376 : entity work.gfmul
port map(
a=>a_2,
b=>"1011010011",
X=>mulr_2_376);

mulc_3_376 : entity work.gfmul
port map(
a=>a_3,
b=>"0010100011",
X=>mulr_3_376);

mulc_4_376 : entity work.gfmul
port map(
a=>a_4,
b=>"1010110000",
X=>mulr_4_376);

mulr_1_377<=a_1;
mulc_2_377 : entity work.gfmul
port map(
a=>a_2,
b=>"0110101111",
X=>mulr_2_377);

mulc_3_377 : entity work.gfmul
port map(
a=>a_3,
b=>"1010001100",
X=>mulr_3_377);

mulc_4_377 : entity work.gfmul
port map(
a=>a_4,
b=>"0110101101",
X=>mulr_4_377);

mulr_1_378<=a_1;
mulc_2_378 : entity work.gfmul
port map(
a=>a_2,
b=>"1101011110",
X=>mulr_2_378);

mulc_3_378 : entity work.gfmul
port map(
a=>a_3,
b=>"1000100010",
X=>mulr_3_378);

mulc_4_378 : entity work.gfmul
port map(
a=>a_4,
b=>"0101110011",
X=>mulr_4_378);

mulr_1_379<=a_1;
mulc_2_379 : entity work.gfmul
port map(
a=>a_2,
b=>"1010110101",
X=>mulr_2_379);

mulc_3_379 : entity work.gfmul
port map(
a=>a_3,
b=>"0010011010",
X=>mulr_3_379);

mulc_4_379 : entity work.gfmul
port map(
a=>a_4,
b=>"1110001010",
X=>mulr_4_379);

mulr_1_380<=a_1;
mulc_2_380 : entity work.gfmul
port map(
a=>a_2,
b=>"0101100011",
X=>mulr_2_380);

mulc_3_380 : entity work.gfmul
port map(
a=>a_3,
b=>"1001101000",
X=>mulr_3_380);

mulc_4_380 : entity work.gfmul
port map(
a=>a_4,
b=>"0001101111",
X=>mulr_4_380);

mulr_1_381<=a_1;
mulc_2_381 : entity work.gfmul
port map(
a=>a_2,
b=>"1011000110",
X=>mulr_2_381);

mulc_3_381 : entity work.gfmul
port map(
a=>a_3,
b=>"0110110010",
X=>mulr_3_381);

mulc_4_381 : entity work.gfmul
port map(
a=>a_4,
b=>"1101111000",
X=>mulr_4_381);

mulr_1_382<=a_1;
mulc_2_382 : entity work.gfmul
port map(
a=>a_2,
b=>"0110000101",
X=>mulr_2_382);

mulc_3_382 : entity work.gfmul
port map(
a=>a_3,
b=>"1011000001",
X=>mulr_3_382);

mulc_4_382 : entity work.gfmul
port map(
a=>a_4,
b=>"1111110110",
X=>mulr_4_382);

mulr_1_383<=a_1;
mulc_2_383 : entity work.gfmul
port map(
a=>a_2,
b=>"1100001010",
X=>mulr_2_383);

mulc_3_383 : entity work.gfmul
port map(
a=>a_3,
b=>"1100010110",
X=>mulr_3_383);

mulc_4_383 : entity work.gfmul
port map(
a=>a_4,
b=>"1110001111",
X=>mulr_4_383);

mulr_1_384<=a_1;
mulc_2_384 : entity work.gfmul
port map(
a=>a_2,
b=>"1000011101",
X=>mulr_2_384);

mulc_3_384 : entity work.gfmul
port map(
a=>a_3,
b=>"0001000011",
X=>mulr_3_384);

mulc_4_384 : entity work.gfmul
port map(
a=>a_4,
b=>"0001000111",
X=>mulr_4_384);

mulr_1_385<=a_1;
mulc_2_385 : entity work.gfmul
port map(
a=>a_2,
b=>"0000110011",
X=>mulr_2_385);

mulc_3_385 : entity work.gfmul
port map(
a=>a_3,
b=>"0100001100",
X=>mulr_3_385);

mulc_4_385 : entity work.gfmul
port map(
a=>a_4,
b=>"1000111000",
X=>mulr_4_385);

mulr_1_386<=a_1;
mulc_2_386 : entity work.gfmul
port map(
a=>a_2,
b=>"0001100110",
X=>mulr_2_386);

mulc_3_386 : entity work.gfmul
port map(
a=>a_3,
b=>"0000111001",
X=>mulr_3_386);

mulc_4_386 : entity work.gfmul
port map(
a=>a_4,
b=>"0111100100",
X=>mulr_4_386);

mulr_1_387<=a_1;
mulc_2_387 : entity work.gfmul
port map(
a=>a_2,
b=>"0011001100",
X=>mulr_2_387);

mulc_3_387 : entity work.gfmul
port map(
a=>a_3,
b=>"0011100100",
X=>mulr_3_387);

mulc_4_387 : entity work.gfmul
port map(
a=>a_4,
b=>"1100111011",
X=>mulr_4_387);

mulr_1_388<=a_1;
mulc_2_388 : entity work.gfmul
port map(
a=>a_2,
b=>"0110011000",
X=>mulr_2_388);

mulc_3_388 : entity work.gfmul
port map(
a=>a_3,
b=>"1110010000",
X=>mulr_3_388);

mulc_4_388 : entity work.gfmul
port map(
a=>a_4,
b=>"0111101110",
X=>mulr_4_388);

mulr_1_389<=a_1;
mulc_2_389 : entity work.gfmul
port map(
a=>a_2,
b=>"1100110000",
X=>mulr_2_389);

mulc_3_389 : entity work.gfmul
port map(
a=>a_3,
b=>"1001011011",
X=>mulr_3_389);

mulc_4_389 : entity work.gfmul
port map(
a=>a_4,
b=>"1101101011",
X=>mulr_4_389);

mulr_1_390<=a_1;
mulc_2_390 : entity work.gfmul
port map(
a=>a_2,
b=>"1001101001",
X=>mulr_2_390);

mulc_3_390 : entity work.gfmul
port map(
a=>a_3,
b=>"0101111110",
X=>mulr_3_390);

mulc_4_390 : entity work.gfmul
port map(
a=>a_4,
b=>"1101101110",
X=>mulr_4_390);

mulr_1_391<=a_1;
mulc_2_391 : entity work.gfmul
port map(
a=>a_2,
b=>"0011011011",
X=>mulr_2_391);

mulc_3_391 : entity work.gfmul
port map(
a=>a_3,
b=>"0111110001",
X=>mulr_3_391);

mulc_4_391 : entity work.gfmul
port map(
a=>a_4,
b=>"1101000110",
X=>mulr_4_391);

mulr_1_392<=a_1;
mulc_2_392 : entity work.gfmul
port map(
a=>a_2,
b=>"0110110110",
X=>mulr_2_392);

mulc_3_392 : entity work.gfmul
port map(
a=>a_3,
b=>"1111001101",
X=>mulr_3_392);

mulc_4_392 : entity work.gfmul
port map(
a=>a_4,
b=>"1000000110",
X=>mulr_4_392);

mulr_1_393<=a_1;
mulc_2_393 : entity work.gfmul
port map(
a=>a_2,
b=>"1101101100",
X=>mulr_2_393);

mulc_3_393 : entity work.gfmul
port map(
a=>a_3,
b=>"1100101111",
X=>mulr_3_393);

mulc_4_393 : entity work.gfmul
port map(
a=>a_4,
b=>"0000010100",
X=>mulr_4_393);

mulr_1_394<=a_1;
mulc_2_394 : entity work.gfmul
port map(
a=>a_2,
b=>"1011010001",
X=>mulr_2_394);

mulc_3_394 : entity work.gfmul
port map(
a=>a_3,
b=>"0010100111",
X=>mulr_3_394);

mulc_4_394 : entity work.gfmul
port map(
a=>a_4,
b=>"0010100000",
X=>mulr_4_394);

mulr_1_395<=a_1;
mulc_2_395 : entity work.gfmul
port map(
a=>a_2,
b=>"0110101011",
X=>mulr_2_395);

mulc_3_395 : entity work.gfmul
port map(
a=>a_3,
b=>"1010011100",
X=>mulr_3_395);

mulc_4_395 : entity work.gfmul
port map(
a=>a_4,
b=>"0100001001",
X=>mulr_4_395);

mulr_1_396<=a_1;
mulc_2_396 : entity work.gfmul
port map(
a=>a_2,
b=>"1101010110",
X=>mulr_2_396);

mulc_3_396 : entity work.gfmul
port map(
a=>a_3,
b=>"1001100010",
X=>mulr_3_396);

mulc_4_396 : entity work.gfmul
port map(
a=>a_4,
b=>"0001011010",
X=>mulr_4_396);

mulr_1_397<=a_1;
mulc_2_397 : entity work.gfmul
port map(
a=>a_2,
b=>"1010100101",
X=>mulr_2_397);

mulc_3_397 : entity work.gfmul
port map(
a=>a_3,
b=>"0110011010",
X=>mulr_3_397);

mulc_4_397 : entity work.gfmul
port map(
a=>a_4,
b=>"1011010000",
X=>mulr_4_397);

mulr_1_398<=a_1;
mulc_2_398 : entity work.gfmul
port map(
a=>a_2,
b=>"0101000011",
X=>mulr_2_398);

mulc_3_398 : entity work.gfmul
port map(
a=>a_3,
b=>"1001100001",
X=>mulr_3_398);

mulc_4_398 : entity work.gfmul
port map(
a=>a_4,
b=>"1010101101",
X=>mulr_4_398);

mulr_1_399<=a_1;
mulc_2_399 : entity work.gfmul
port map(
a=>a_2,
b=>"1010000110",
X=>mulr_2_399);

mulc_3_399 : entity work.gfmul
port map(
a=>a_3,
b=>"0110010110",
X=>mulr_3_399);

mulc_4_399 : entity work.gfmul
port map(
a=>a_4,
b=>"0101000101",
X=>mulr_4_399);

mulr_1_400<=a_1;
mulc_2_400 : entity work.gfmul
port map(
a=>a_2,
b=>"0100000101",
X=>mulr_2_400);

mulc_3_400 : entity work.gfmul
port map(
a=>a_3,
b=>"1001010001",
X=>mulr_3_400);

mulc_4_400 : entity work.gfmul
port map(
a=>a_4,
b=>"1000111010",
X=>mulr_4_400);

mulr_1_401<=a_1;
mulc_2_401 : entity work.gfmul
port map(
a=>a_2,
b=>"1000001010",
X=>mulr_2_401);

mulc_3_401 : entity work.gfmul
port map(
a=>a_3,
b=>"0101010110",
X=>mulr_3_401);

mulc_4_401 : entity work.gfmul
port map(
a=>a_4,
b=>"0111110100",
X=>mulr_4_401);

mulr_1_402<=a_1;
mulc_2_402 : entity work.gfmul
port map(
a=>a_2,
b=>"0000011101",
X=>mulr_2_402);

mulc_3_402 : entity work.gfmul
port map(
a=>a_3,
b=>"0101010001",
X=>mulr_3_402);

mulc_4_402 : entity work.gfmul
port map(
a=>a_4,
b=>"1110111011",
X=>mulr_4_402);

mulr_1_403<=a_1;
mulc_2_403 : entity work.gfmul
port map(
a=>a_2,
b=>"0000111010",
X=>mulr_2_403);

mulc_3_403 : entity work.gfmul
port map(
a=>a_3,
b=>"0101001101",
X=>mulr_3_403);

mulc_4_403 : entity work.gfmul
port map(
a=>a_4,
b=>"0111100111",
X=>mulr_4_403);

mulr_1_404<=a_1;
mulc_2_404 : entity work.gfmul
port map(
a=>a_2,
b=>"0001110100",
X=>mulr_2_404);

mulc_3_404 : entity work.gfmul
port map(
a=>a_3,
b=>"0100111101",
X=>mulr_3_404);

mulc_4_404 : entity work.gfmul
port map(
a=>a_4,
b=>"1100100011",
X=>mulr_4_404);

mulr_1_405<=a_1;
mulc_2_405 : entity work.gfmul
port map(
a=>a_2,
b=>"0011101000",
X=>mulr_2_405);

mulc_3_405 : entity work.gfmul
port map(
a=>a_3,
b=>"0011111101",
X=>mulr_3_405);

mulc_4_405 : entity work.gfmul
port map(
a=>a_4,
b=>"0100101110",
X=>mulr_4_405);

mulr_1_406<=a_1;
mulc_2_406 : entity work.gfmul
port map(
a=>a_2,
b=>"0111010000",
X=>mulr_2_406);

mulc_3_406 : entity work.gfmul
port map(
a=>a_3,
b=>"1111110100",
X=>mulr_3_406);

mulc_4_406 : entity work.gfmul
port map(
a=>a_4,
b=>"0101100010",
X=>mulr_4_406);

mulr_1_407<=a_1;
mulc_2_407 : entity work.gfmul
port map(
a=>a_2,
b=>"1110100000",
X=>mulr_2_407);

mulc_3_407 : entity work.gfmul
port map(
a=>a_3,
b=>"1111001011",
X=>mulr_3_407);

mulc_4_407 : entity work.gfmul
port map(
a=>a_4,
b=>"1100000010",
X=>mulr_4_407);

mulr_1_408<=a_1;
mulc_2_408 : entity work.gfmul
port map(
a=>a_2,
b=>"1101001001",
X=>mulr_2_408);

mulc_3_408 : entity work.gfmul
port map(
a=>a_3,
b=>"1100110111",
X=>mulr_3_408);

mulc_4_408 : entity work.gfmul
port map(
a=>a_4,
b=>"0000100110",
X=>mulr_4_408);

mulr_1_409<=a_1;
mulc_2_409 : entity work.gfmul
port map(
a=>a_2,
b=>"1010011011",
X=>mulr_2_409);

mulc_3_409 : entity work.gfmul
port map(
a=>a_3,
b=>"0011000111",
X=>mulr_3_409);

mulc_4_409 : entity work.gfmul
port map(
a=>a_4,
b=>"0100110000",
X=>mulr_4_409);

mulr_1_410<=a_1;
mulc_2_410 : entity work.gfmul
port map(
a=>a_2,
b=>"0100111111",
X=>mulr_2_410);

mulc_3_410 : entity work.gfmul
port map(
a=>a_3,
b=>"1100011100",
X=>mulr_3_410);

mulc_4_410 : entity work.gfmul
port map(
a=>a_4,
b=>"0110010010",
X=>mulr_4_410);

mulr_1_411<=a_1;
mulc_2_411 : entity work.gfmul
port map(
a=>a_2,
b=>"1001111110",
X=>mulr_2_411);

mulc_3_411 : entity work.gfmul
port map(
a=>a_3,
b=>"0001101011",
X=>mulr_3_411);

mulc_4_411 : entity work.gfmul
port map(
a=>a_4,
b=>"0010001011",
X=>mulr_4_411);

mulr_1_412<=a_1;
mulc_2_412 : entity work.gfmul
port map(
a=>a_2,
b=>"0011110101",
X=>mulr_2_412);

mulc_3_412 : entity work.gfmul
port map(
a=>a_3,
b=>"0110101100",
X=>mulr_3_412);

mulc_4_412 : entity work.gfmul
port map(
a=>a_4,
b=>"0001010001",
X=>mulr_4_412);

mulr_1_413<=a_1;
mulc_2_413 : entity work.gfmul
port map(
a=>a_2,
b=>"0111101010",
X=>mulr_2_413);

mulc_3_413 : entity work.gfmul
port map(
a=>a_3,
b=>"1010111001",
X=>mulr_3_413);

mulc_4_413 : entity work.gfmul
port map(
a=>a_4,
b=>"1010001000",
X=>mulr_4_413);

mulr_1_414<=a_1;
mulc_2_414 : entity work.gfmul
port map(
a=>a_2,
b=>"1111010100",
X=>mulr_2_414);

mulc_3_414 : entity work.gfmul
port map(
a=>a_3,
b=>"1011110110",
X=>mulr_3_414);

mulc_4_414 : entity work.gfmul
port map(
a=>a_4,
b=>"0001101101",
X=>mulr_4_414);

mulr_1_415<=a_1;
mulc_2_415 : entity work.gfmul
port map(
a=>a_2,
b=>"1110100001",
X=>mulr_2_415);

mulc_3_415 : entity work.gfmul
port map(
a=>a_3,
b=>"1111001010",
X=>mulr_3_415);

mulc_4_415 : entity work.gfmul
port map(
a=>a_4,
b=>"1101101000",
X=>mulr_4_415);

mulr_1_416<=a_1;
mulc_2_416 : entity work.gfmul
port map(
a=>a_2,
b=>"1101001011",
X=>mulr_2_416);

mulc_3_416 : entity work.gfmul
port map(
a=>a_3,
b=>"1100110011",
X=>mulr_3_416);

mulc_4_416 : entity work.gfmul
port map(
a=>a_4,
b=>"1101110110",
X=>mulr_4_416);

mulr_1_417<=a_1;
mulc_2_417 : entity work.gfmul
port map(
a=>a_2,
b=>"1010011111",
X=>mulr_2_417);

mulc_3_417 : entity work.gfmul
port map(
a=>a_3,
b=>"0011010111",
X=>mulr_3_417);

mulc_4_417 : entity work.gfmul
port map(
a=>a_4,
b=>"1110000110",
X=>mulr_4_417);

mulr_1_418<=a_1;
mulc_2_418 : entity work.gfmul
port map(
a=>a_2,
b=>"0100110111",
X=>mulr_2_418);

mulc_3_418 : entity work.gfmul
port map(
a=>a_3,
b=>"1101011100",
X=>mulr_3_418);

mulc_4_418 : entity work.gfmul
port map(
a=>a_4,
b=>"0000001111",
X=>mulr_4_418);

mulr_1_419<=a_1;
mulc_2_419 : entity work.gfmul
port map(
a=>a_2,
b=>"1001101110",
X=>mulr_2_419);

mulc_3_419 : entity work.gfmul
port map(
a=>a_3,
b=>"0101101011",
X=>mulr_3_419);

mulc_4_419 : entity work.gfmul
port map(
a=>a_4,
b=>"0001111000",
X=>mulr_4_419);

mulr_1_420<=a_1;
mulc_2_420 : entity work.gfmul
port map(
a=>a_2,
b=>"0011010101",
X=>mulr_2_420);

mulc_3_420 : entity work.gfmul
port map(
a=>a_3,
b=>"0110100101",
X=>mulr_3_420);

mulc_4_420 : entity work.gfmul
port map(
a=>a_4,
b=>"1111000000",
X=>mulr_4_420);

mulr_1_421<=a_1;
mulc_2_421 : entity work.gfmul
port map(
a=>a_2,
b=>"0110101010",
X=>mulr_2_421);

mulc_3_421 : entity work.gfmul
port map(
a=>a_3,
b=>"1010011101",
X=>mulr_3_421);

mulc_4_421 : entity work.gfmul
port map(
a=>a_4,
b=>"1000111111",
X=>mulr_4_421);

mulr_1_422<=a_1;
mulc_2_422 : entity work.gfmul
port map(
a=>a_2,
b=>"1101010100",
X=>mulr_2_422);

mulc_3_422 : entity work.gfmul
port map(
a=>a_3,
b=>"1001100110",
X=>mulr_3_422);

mulc_4_422 : entity work.gfmul
port map(
a=>a_4,
b=>"0111011100",
X=>mulr_4_422);

mulr_1_423<=a_1;
mulc_2_423 : entity work.gfmul
port map(
a=>a_2,
b=>"1010100001",
X=>mulr_2_423);

mulc_3_423 : entity work.gfmul
port map(
a=>a_3,
b=>"0110001010",
X=>mulr_3_423);

mulc_4_423 : entity work.gfmul
port map(
a=>a_4,
b=>"1011111011",
X=>mulr_4_423);

mulr_1_424<=a_1;
mulc_2_424 : entity work.gfmul
port map(
a=>a_2,
b=>"0101001011",
X=>mulr_2_424);

mulc_3_424 : entity work.gfmul
port map(
a=>a_3,
b=>"1000100001",
X=>mulr_3_424);

mulc_4_424 : entity work.gfmul
port map(
a=>a_4,
b=>"1111110101",
X=>mulr_4_424);

mulr_1_425<=a_1;
mulc_2_425 : entity work.gfmul
port map(
a=>a_2,
b=>"1010010110",
X=>mulr_2_425);

mulc_3_425 : entity work.gfmul
port map(
a=>a_3,
b=>"0010010110",
X=>mulr_3_425);

mulc_4_425 : entity work.gfmul
port map(
a=>a_4,
b=>"1110010111",
X=>mulr_4_425);

mulr_1_426<=a_1;
mulc_2_426 : entity work.gfmul
port map(
a=>a_2,
b=>"0100100101",
X=>mulr_2_426);

mulc_3_426 : entity work.gfmul
port map(
a=>a_3,
b=>"1001011000",
X=>mulr_3_426);

mulc_4_426 : entity work.gfmul
port map(
a=>a_4,
b=>"0010000111",
X=>mulr_4_426);

mulr_1_427<=a_1;
mulc_2_427 : entity work.gfmul
port map(
a=>a_2,
b=>"1001001010",
X=>mulr_2_427);

mulc_3_427 : entity work.gfmul
port map(
a=>a_3,
b=>"0101110010",
X=>mulr_3_427);

mulc_4_427 : entity work.gfmul
port map(
a=>a_4,
b=>"0000110001",
X=>mulr_4_427);

mulr_1_428<=a_1;
mulc_2_428 : entity work.gfmul
port map(
a=>a_2,
b=>"0010011101",
X=>mulr_2_428);

mulc_3_428 : entity work.gfmul
port map(
a=>a_3,
b=>"0111000001",
X=>mulr_3_428);

mulc_4_428 : entity work.gfmul
port map(
a=>a_4,
b=>"0110001000",
X=>mulr_4_428);

mulr_1_429<=a_1;
mulc_2_429 : entity work.gfmul
port map(
a=>a_2,
b=>"0100111010",
X=>mulr_2_429);

mulc_3_429 : entity work.gfmul
port map(
a=>a_3,
b=>"1100001101",
X=>mulr_3_429);

mulc_4_429 : entity work.gfmul
port map(
a=>a_4,
b=>"0001011011",
X=>mulr_4_429);

mulr_1_430<=a_1;
mulc_2_430 : entity work.gfmul
port map(
a=>a_2,
b=>"1001110100",
X=>mulr_2_430);

mulc_3_430 : entity work.gfmul
port map(
a=>a_3,
b=>"0000101111",
X=>mulr_3_430);

mulc_4_430 : entity work.gfmul
port map(
a=>a_4,
b=>"1011011000",
X=>mulr_4_430);

mulr_1_431<=a_1;
mulc_2_431 : entity work.gfmul
port map(
a=>a_2,
b=>"0011100001",
X=>mulr_2_431);

mulc_3_431 : entity work.gfmul
port map(
a=>a_3,
b=>"0010111100",
X=>mulr_3_431);

mulc_4_431 : entity work.gfmul
port map(
a=>a_4,
b=>"1011101101",
X=>mulr_4_431);

mulr_1_432<=a_1;
mulc_2_432 : entity work.gfmul
port map(
a=>a_2,
b=>"0111000010",
X=>mulr_2_432);

mulc_3_432 : entity work.gfmul
port map(
a=>a_3,
b=>"1011110000",
X=>mulr_3_432);

mulc_4_432 : entity work.gfmul
port map(
a=>a_4,
b=>"1101000101",
X=>mulr_4_432);

mulr_1_433<=a_1;
mulc_2_433 : entity work.gfmul
port map(
a=>a_2,
b=>"1110000100",
X=>mulr_2_433);

mulc_3_433 : entity work.gfmul
port map(
a=>a_3,
b=>"1111010010",
X=>mulr_3_433);

mulc_4_433 : entity work.gfmul
port map(
a=>a_4,
b=>"1000011110",
X=>mulr_4_433);

mulr_1_434<=a_1;
mulc_2_434 : entity work.gfmul
port map(
a=>a_2,
b=>"1100000001",
X=>mulr_2_434);

mulc_3_434 : entity work.gfmul
port map(
a=>a_3,
b=>"1101010011",
X=>mulr_3_434);

mulc_4_434 : entity work.gfmul
port map(
a=>a_4,
b=>"0011010100",
X=>mulr_4_434);

mulr_1_435<=a_1;
mulc_2_435 : entity work.gfmul
port map(
a=>a_2,
b=>"1000001011",
X=>mulr_2_435);

mulc_3_435 : entity work.gfmul
port map(
a=>a_3,
b=>"0101010111",
X=>mulr_3_435);

mulc_4_435 : entity work.gfmul
port map(
a=>a_4,
b=>"1010101001",
X=>mulr_4_435);

mulr_1_436<=a_1;
mulc_2_436 : entity work.gfmul
port map(
a=>a_2,
b=>"0000011111",
X=>mulr_2_436);

mulc_3_436 : entity work.gfmul
port map(
a=>a_3,
b=>"0101010101",
X=>mulr_3_436);

mulc_4_436 : entity work.gfmul
port map(
a=>a_4,
b=>"0101100101",
X=>mulr_4_436);

mulr_1_437<=a_1;
mulc_2_437 : entity work.gfmul
port map(
a=>a_2,
b=>"0000111110",
X=>mulr_2_437);

mulc_3_437 : entity work.gfmul
port map(
a=>a_3,
b=>"0101011101",
X=>mulr_3_437);

mulc_4_437 : entity work.gfmul
port map(
a=>a_4,
b=>"1100111010",
X=>mulr_4_437);

mulr_1_438<=a_1;
mulc_2_438 : entity work.gfmul
port map(
a=>a_2,
b=>"0001111100",
X=>mulr_2_438);

mulc_3_438 : entity work.gfmul
port map(
a=>a_3,
b=>"0101111101",
X=>mulr_3_438);

mulc_4_438 : entity work.gfmul
port map(
a=>a_4,
b=>"0111100110",
X=>mulr_4_438);

mulr_1_439<=a_1;
mulc_2_439 : entity work.gfmul
port map(
a=>a_2,
b=>"0011111000",
X=>mulr_2_439);

mulc_3_439 : entity work.gfmul
port map(
a=>a_3,
b=>"0111111101",
X=>mulr_3_439);

mulc_4_439 : entity work.gfmul
port map(
a=>a_4,
b=>"1100101011",
X=>mulr_4_439);

mulr_1_440<=a_1;
mulc_2_440 : entity work.gfmul
port map(
a=>a_2,
b=>"0111110000",
X=>mulr_2_440);

mulc_3_440 : entity work.gfmul
port map(
a=>a_3,
b=>"1111111101",
X=>mulr_3_440);

mulc_4_440 : entity work.gfmul
port map(
a=>a_4,
b=>"0101101110",
X=>mulr_4_440);

mulr_1_441<=a_1;
mulc_2_441 : entity work.gfmul
port map(
a=>a_2,
b=>"1111100000",
X=>mulr_2_441);

mulc_3_441 : entity work.gfmul
port map(
a=>a_3,
b=>"1111101111",
X=>mulr_3_441);

mulc_4_441 : entity work.gfmul
port map(
a=>a_4,
b=>"1101100010",
X=>mulr_4_441);

mulr_1_442<=a_1;
mulc_2_442 : entity work.gfmul
port map(
a=>a_2,
b=>"1111001001",
X=>mulr_2_442);

mulc_3_442 : entity work.gfmul
port map(
a=>a_3,
b=>"1110100111",
X=>mulr_3_442);

mulc_4_442 : entity work.gfmul
port map(
a=>a_4,
b=>"1100100110",
X=>mulr_4_442);

mulr_1_443<=a_1;
mulc_2_443 : entity work.gfmul
port map(
a=>a_2,
b=>"1110011011",
X=>mulr_2_443);

mulc_3_443 : entity work.gfmul
port map(
a=>a_3,
b=>"1010000111",
X=>mulr_3_443);

mulc_4_443 : entity work.gfmul
port map(
a=>a_4,
b=>"0100000110",
X=>mulr_4_443);

mulr_1_444<=a_1;
mulc_2_444 : entity work.gfmul
port map(
a=>a_2,
b=>"1100111111",
X=>mulr_2_444);

mulc_3_444 : entity work.gfmul
port map(
a=>a_3,
b=>"1000001110",
X=>mulr_3_444);

mulc_4_444 : entity work.gfmul
port map(
a=>a_4,
b=>"0000100010",
X=>mulr_4_444);

mulr_1_445<=a_1;
mulc_2_445 : entity work.gfmul
port map(
a=>a_2,
b=>"1001110111",
X=>mulr_2_445);

mulc_3_445 : entity work.gfmul
port map(
a=>a_3,
b=>"0000101010",
X=>mulr_3_445);

mulc_4_445 : entity work.gfmul
port map(
a=>a_4,
b=>"0100010000",
X=>mulr_4_445);

mulr_1_446<=a_1;
mulc_2_446 : entity work.gfmul
port map(
a=>a_2,
b=>"0011100111",
X=>mulr_2_446);

mulc_3_446 : entity work.gfmul
port map(
a=>a_3,
b=>"0010101000",
X=>mulr_3_446);

mulc_4_446 : entity work.gfmul
port map(
a=>a_4,
b=>"0010010010",
X=>mulr_4_446);

mulr_1_447<=a_1;
mulc_2_447 : entity work.gfmul
port map(
a=>a_2,
b=>"0111001110",
X=>mulr_2_447);

mulc_3_447 : entity work.gfmul
port map(
a=>a_3,
b=>"1010100000",
X=>mulr_3_447);

mulc_4_447 : entity work.gfmul
port map(
a=>a_4,
b=>"0010011001",
X=>mulr_4_447);

mulr_1_448<=a_1;
mulc_2_448 : entity work.gfmul
port map(
a=>a_2,
b=>"1110011100",
X=>mulr_2_448);

mulc_3_448 : entity work.gfmul
port map(
a=>a_3,
b=>"1010010010",
X=>mulr_3_448);

mulc_4_448 : entity work.gfmul
port map(
a=>a_4,
b=>"0011000001",
X=>mulr_4_448);

mulr_1_449<=a_1;
mulc_2_449 : entity work.gfmul
port map(
a=>a_2,
b=>"1100110001",
X=>mulr_2_449);

mulc_3_449 : entity work.gfmul
port map(
a=>a_3,
b=>"1001011010",
X=>mulr_3_449);

mulc_4_449 : entity work.gfmul
port map(
a=>a_4,
b=>"1000000001",
X=>mulr_4_449);

mulr_1_450<=a_1;
mulc_2_450 : entity work.gfmul
port map(
a=>a_2,
b=>"1001101011",
X=>mulr_2_450);

mulc_3_450 : entity work.gfmul
port map(
a=>a_3,
b=>"0101111010",
X=>mulr_3_450);

mulc_4_450 : entity work.gfmul
port map(
a=>a_4,
b=>"0000101100",
X=>mulr_4_450);

mulr_1_451<=a_1;
mulc_2_451 : entity work.gfmul
port map(
a=>a_2,
b=>"0011011111",
X=>mulr_2_451);

mulc_3_451 : entity work.gfmul
port map(
a=>a_3,
b=>"0111100001",
X=>mulr_3_451);

mulc_4_451 : entity work.gfmul
port map(
a=>a_4,
b=>"0101100000",
X=>mulr_4_451);

mulr_1_452<=a_1;
mulc_2_452 : entity work.gfmul
port map(
a=>a_2,
b=>"0110111110",
X=>mulr_2_452);

mulc_3_452 : entity work.gfmul
port map(
a=>a_3,
b=>"1110001101",
X=>mulr_3_452);

mulc_4_452 : entity work.gfmul
port map(
a=>a_4,
b=>"1100010010",
X=>mulr_4_452);

mulr_1_453<=a_1;
mulc_2_453 : entity work.gfmul
port map(
a=>a_2,
b=>"1101111100",
X=>mulr_2_453);

mulc_3_453 : entity work.gfmul
port map(
a=>a_3,
b=>"1000101111",
X=>mulr_3_453);

mulc_4_453 : entity work.gfmul
port map(
a=>a_4,
b=>"0010100110",
X=>mulr_4_453);

mulr_1_454<=a_1;
mulc_2_454 : entity work.gfmul
port map(
a=>a_2,
b=>"1011110001",
X=>mulr_2_454);

mulc_3_454 : entity work.gfmul
port map(
a=>a_3,
b=>"0010101110",
X=>mulr_3_454);

mulc_4_454 : entity work.gfmul
port map(
a=>a_4,
b=>"0100111001",
X=>mulr_4_454);

mulr_1_455<=a_1;
mulc_2_455 : entity work.gfmul
port map(
a=>a_2,
b=>"0111101011",
X=>mulr_2_455);

mulc_3_455 : entity work.gfmul
port map(
a=>a_3,
b=>"1010111000",
X=>mulr_3_455);

mulc_4_455 : entity work.gfmul
port map(
a=>a_4,
b=>"0111011010",
X=>mulr_4_455);

mulr_1_456<=a_1;
mulc_2_456 : entity work.gfmul
port map(
a=>a_2,
b=>"1111010110",
X=>mulr_2_456);

mulc_3_456 : entity work.gfmul
port map(
a=>a_3,
b=>"1011110010",
X=>mulr_3_456);

mulc_4_456 : entity work.gfmul
port map(
a=>a_4,
b=>"1011001011",
X=>mulr_4_456);

mulr_1_457<=a_1;
mulc_2_457 : entity work.gfmul
port map(
a=>a_2,
b=>"1110100101",
X=>mulr_2_457);

mulc_3_457 : entity work.gfmul
port map(
a=>a_3,
b=>"1111011010",
X=>mulr_3_457);

mulc_4_457 : entity work.gfmul
port map(
a=>a_4,
b=>"1001110101",
X=>mulr_4_457);

mulr_1_458<=a_1;
mulc_2_458 : entity work.gfmul
port map(
a=>a_2,
b=>"1101000011",
X=>mulr_2_458);

mulc_3_458 : entity work.gfmul
port map(
a=>a_3,
b=>"1101110011",
X=>mulr_3_458);

mulc_4_458 : entity work.gfmul
port map(
a=>a_4,
b=>"1110001100",
X=>mulr_4_458);

mulr_1_459<=a_1;
mulc_2_459 : entity work.gfmul
port map(
a=>a_2,
b=>"1010001111",
X=>mulr_2_459);

mulc_3_459 : entity work.gfmul
port map(
a=>a_3,
b=>"0111010111",
X=>mulr_3_459);

mulc_4_459 : entity work.gfmul
port map(
a=>a_4,
b=>"0001011111",
X=>mulr_4_459);

mulr_1_460<=a_1;
mulc_2_460 : entity work.gfmul
port map(
a=>a_2,
b=>"0100010111",
X=>mulr_2_460);

mulc_3_460 : entity work.gfmul
port map(
a=>a_3,
b=>"1101010101",
X=>mulr_3_460);

mulc_4_460 : entity work.gfmul
port map(
a=>a_4,
b=>"1011111000",
X=>mulr_4_460);

mulr_1_461<=a_1;
mulc_2_461 : entity work.gfmul
port map(
a=>a_2,
b=>"1000101110",
X=>mulr_2_461);

mulc_3_461 : entity work.gfmul
port map(
a=>a_3,
b=>"0101001111",
X=>mulr_3_461);

mulc_4_461 : entity work.gfmul
port map(
a=>a_4,
b=>"1111101101",
X=>mulr_4_461);

mulr_1_462<=a_1;
mulc_2_462 : entity work.gfmul
port map(
a=>a_2,
b=>"0001010101",
X=>mulr_2_462);

mulc_3_462 : entity work.gfmul
port map(
a=>a_3,
b=>"0100110101",
X=>mulr_3_462);

mulc_4_462 : entity work.gfmul
port map(
a=>a_4,
b=>"1101010111",
X=>mulr_4_462);

mulr_1_463<=a_1;
mulc_2_463 : entity work.gfmul
port map(
a=>a_2,
b=>"0010101010",
X=>mulr_2_463);

mulc_3_463 : entity work.gfmul
port map(
a=>a_3,
b=>"0011011101",
X=>mulr_3_463);

mulc_4_463 : entity work.gfmul
port map(
a=>a_4,
b=>"1010001110",
X=>mulr_4_463);

mulr_1_464<=a_1;
mulc_2_464 : entity work.gfmul
port map(
a=>a_2,
b=>"0101010100",
X=>mulr_2_464);

mulc_3_464 : entity work.gfmul
port map(
a=>a_3,
b=>"1101110100",
X=>mulr_3_464);

mulc_4_464 : entity work.gfmul
port map(
a=>a_4,
b=>"0001011101",
X=>mulr_4_464);

mulr_1_465<=a_1;
mulc_2_465 : entity work.gfmul
port map(
a=>a_2,
b=>"1010101000",
X=>mulr_2_465);

mulc_3_465 : entity work.gfmul
port map(
a=>a_3,
b=>"0111001011",
X=>mulr_3_465);

mulc_4_465 : entity work.gfmul
port map(
a=>a_4,
b=>"1011101000",
X=>mulr_4_465);

mulr_1_466<=a_1;
mulc_2_466 : entity work.gfmul
port map(
a=>a_2,
b=>"0101011001",
X=>mulr_2_466);

mulc_3_466 : entity work.gfmul
port map(
a=>a_3,
b=>"1100100101",
X=>mulr_3_466);

mulc_4_466 : entity work.gfmul
port map(
a=>a_4,
b=>"1101101101",
X=>mulr_4_466);

mulr_1_467<=a_1;
mulc_2_467 : entity work.gfmul
port map(
a=>a_2,
b=>"1010110010",
X=>mulr_2_467);

mulc_3_467 : entity work.gfmul
port map(
a=>a_3,
b=>"0010001111",
X=>mulr_3_467);

mulc_4_467 : entity work.gfmul
port map(
a=>a_4,
b=>"1101011110",
X=>mulr_4_467);

mulr_1_468<=a_1;
mulc_2_468 : entity work.gfmul
port map(
a=>a_2,
b=>"0101101101",
X=>mulr_2_468);

mulc_3_468 : entity work.gfmul
port map(
a=>a_3,
b=>"1000111100",
X=>mulr_3_468);

mulc_4_468 : entity work.gfmul
port map(
a=>a_4,
b=>"1011000110",
X=>mulr_4_468);

mulr_1_469<=a_1;
mulc_2_469 : entity work.gfmul
port map(
a=>a_2,
b=>"1011011010",
X=>mulr_2_469);

mulc_3_469 : entity work.gfmul
port map(
a=>a_3,
b=>"0011100010",
X=>mulr_3_469);

mulc_4_469 : entity work.gfmul
port map(
a=>a_4,
b=>"1000011101",
X=>mulr_4_469);

mulr_1_470<=a_1;
mulc_2_470 : entity work.gfmul
port map(
a=>a_2,
b=>"0110111101",
X=>mulr_2_470);

mulc_3_470 : entity work.gfmul
port map(
a=>a_3,
b=>"1110001000",
X=>mulr_3_470);

mulc_4_470 : entity work.gfmul
port map(
a=>a_4,
b=>"0011001100",
X=>mulr_4_470);

mulr_1_471<=a_1;
mulc_2_471 : entity work.gfmul
port map(
a=>a_2,
b=>"1101111010",
X=>mulr_2_471);

mulc_3_471 : entity work.gfmul
port map(
a=>a_3,
b=>"1000111011",
X=>mulr_3_471);

mulc_4_471 : entity work.gfmul
port map(
a=>a_4,
b=>"1001101001",
X=>mulr_4_471);

mulr_1_472<=a_1;
mulc_2_472 : entity work.gfmul
port map(
a=>a_2,
b=>"1011111101",
X=>mulr_2_472);

mulc_3_472 : entity work.gfmul
port map(
a=>a_3,
b=>"0011111110",
X=>mulr_3_472);

mulc_4_472 : entity work.gfmul
port map(
a=>a_4,
b=>"1101101100",
X=>mulr_4_472);

mulr_1_473<=a_1;
mulc_2_473 : entity work.gfmul
port map(
a=>a_2,
b=>"0111110011",
X=>mulr_2_473);

mulc_3_473 : entity work.gfmul
port map(
a=>a_3,
b=>"1111111000",
X=>mulr_3_473);

mulc_4_473 : entity work.gfmul
port map(
a=>a_4,
b=>"1101010110",
X=>mulr_4_473);

mulr_1_474<=a_1;
mulc_2_474 : entity work.gfmul
port map(
a=>a_2,
b=>"1111100110",
X=>mulr_2_474);

mulc_3_474 : entity work.gfmul
port map(
a=>a_3,
b=>"1111111011",
X=>mulr_3_474);

mulc_4_474 : entity work.gfmul
port map(
a=>a_4,
b=>"1010000110",
X=>mulr_4_474);

mulr_1_475<=a_1;
mulc_2_475 : entity work.gfmul
port map(
a=>a_2,
b=>"1111000101",
X=>mulr_2_475);

mulc_3_475 : entity work.gfmul
port map(
a=>a_3,
b=>"1111110111",
X=>mulr_3_475);

mulc_4_475 : entity work.gfmul
port map(
a=>a_4,
b=>"0000011101",
X=>mulr_4_475);

mulr_1_476<=a_1;
mulc_2_476 : entity work.gfmul
port map(
a=>a_2,
b=>"1110000011",
X=>mulr_2_476);

mulc_3_476 : entity work.gfmul
port map(
a=>a_3,
b=>"1111000111",
X=>mulr_3_476);

mulc_4_476 : entity work.gfmul
port map(
a=>a_4,
b=>"0011101000",
X=>mulr_4_476);

mulr_1_477<=a_1;
mulc_2_477 : entity work.gfmul
port map(
a=>a_2,
b=>"1100001111",
X=>mulr_2_477);

mulc_3_477 : entity work.gfmul
port map(
a=>a_3,
b=>"1100000111",
X=>mulr_3_477);

mulc_4_477 : entity work.gfmul
port map(
a=>a_4,
b=>"1101001001",
X=>mulr_4_477);

mulr_1_478<=a_1;
mulc_2_478 : entity work.gfmul
port map(
a=>a_2,
b=>"1000010111",
X=>mulr_2_478);

mulc_3_478 : entity work.gfmul
port map(
a=>a_3,
b=>"0000000111",
X=>mulr_3_478);

mulc_4_478 : entity work.gfmul
port map(
a=>a_4,
b=>"1001111110",
X=>mulr_4_478);

mulr_1_479<=a_1;
mulc_2_479 : entity work.gfmul
port map(
a=>a_2,
b=>"0000100111",
X=>mulr_2_479);

mulc_3_479 : entity work.gfmul
port map(
a=>a_3,
b=>"0000011100",
X=>mulr_3_479);

mulc_4_479 : entity work.gfmul
port map(
a=>a_4,
b=>"1111010100",
X=>mulr_4_479);

mulr_1_480<=a_1;
mulc_2_480 : entity work.gfmul
port map(
a=>a_2,
b=>"0001001110",
X=>mulr_2_480);

mulc_3_480 : entity work.gfmul
port map(
a=>a_3,
b=>"0001110000",
X=>mulr_3_480);

mulc_4_480 : entity work.gfmul
port map(
a=>a_4,
b=>"1010011111",
X=>mulr_4_480);

mulr_1_481<=a_1;
mulc_2_481 : entity work.gfmul
port map(
a=>a_2,
b=>"0010011100",
X=>mulr_2_481);

mulc_3_481 : entity work.gfmul
port map(
a=>a_3,
b=>"0111000000",
X=>mulr_3_481);

mulc_4_481 : entity work.gfmul
port map(
a=>a_4,
b=>"0011010101",
X=>mulr_4_481);

mulr_1_482<=a_1;
mulc_2_482 : entity work.gfmul
port map(
a=>a_2,
b=>"0100111000",
X=>mulr_2_482);

mulc_3_482 : entity work.gfmul
port map(
a=>a_3,
b=>"1100001001",
X=>mulr_3_482);

mulc_4_482 : entity work.gfmul
port map(
a=>a_4,
b=>"1010100001",
X=>mulr_4_482);

mulr_1_483<=a_1;
mulc_2_483 : entity work.gfmul
port map(
a=>a_2,
b=>"1001110000",
X=>mulr_2_483);

mulc_3_483 : entity work.gfmul
port map(
a=>a_3,
b=>"0000111111",
X=>mulr_3_483);

mulc_4_483 : entity work.gfmul
port map(
a=>a_4,
b=>"0100100101",
X=>mulr_4_483);

mulr_1_484<=a_1;
mulc_2_484 : entity work.gfmul
port map(
a=>a_2,
b=>"0011101001",
X=>mulr_2_484);

mulc_3_484 : entity work.gfmul
port map(
a=>a_3,
b=>"0011111100",
X=>mulr_3_484);

mulc_4_484 : entity work.gfmul
port map(
a=>a_4,
b=>"0100111010",
X=>mulr_4_484);

mulr_1_485<=a_1;
mulc_2_485 : entity work.gfmul
port map(
a=>a_2,
b=>"0111010010",
X=>mulr_2_485);

mulc_3_485 : entity work.gfmul
port map(
a=>a_3,
b=>"1111110000",
X=>mulr_3_485);

mulc_4_485 : entity work.gfmul
port map(
a=>a_4,
b=>"0111000010",
X=>mulr_4_485);

mulr_1_486<=a_1;
mulc_2_486 : entity work.gfmul
port map(
a=>a_2,
b=>"1110100100",
X=>mulr_2_486);

mulc_3_486 : entity work.gfmul
port map(
a=>a_3,
b=>"1111011011",
X=>mulr_3_486);

mulc_4_486 : entity work.gfmul
port map(
a=>a_4,
b=>"1000001011",
X=>mulr_4_486);

mulr_1_487<=a_1;
mulc_2_487 : entity work.gfmul
port map(
a=>a_2,
b=>"1101000001",
X=>mulr_2_487);

mulc_3_487 : entity work.gfmul
port map(
a=>a_3,
b=>"1101110111",
X=>mulr_3_487);

mulc_4_487 : entity work.gfmul
port map(
a=>a_4,
b=>"0001111100",
X=>mulr_4_487);

mulr_1_488<=a_1;
mulc_2_488 : entity work.gfmul
port map(
a=>a_2,
b=>"1010001011",
X=>mulr_2_488);

mulc_3_488 : entity work.gfmul
port map(
a=>a_3,
b=>"0111000111",
X=>mulr_3_488);

mulc_4_488 : entity work.gfmul
port map(
a=>a_4,
b=>"1111100000",
X=>mulr_4_488);

mulr_1_489<=a_1;
mulc_2_489 : entity work.gfmul
port map(
a=>a_2,
b=>"0100011111",
X=>mulr_2_489);

mulc_3_489 : entity work.gfmul
port map(
a=>a_3,
b=>"1100010101",
X=>mulr_3_489);

mulc_4_489 : entity work.gfmul
port map(
a=>a_4,
b=>"1100111111",
X=>mulr_4_489);

mulr_1_490<=a_1;
mulc_2_490 : entity work.gfmul
port map(
a=>a_2,
b=>"1000111110",
X=>mulr_2_490);

mulc_3_490 : entity work.gfmul
port map(
a=>a_3,
b=>"0001001111",
X=>mulr_3_490);

mulc_4_490 : entity work.gfmul
port map(
a=>a_4,
b=>"0111001110",
X=>mulr_4_490);

mulr_1_491<=a_1;
mulc_2_491 : entity work.gfmul
port map(
a=>a_2,
b=>"0001110101",
X=>mulr_2_491);

mulc_3_491 : entity work.gfmul
port map(
a=>a_3,
b=>"0100111100",
X=>mulr_3_491);

mulc_4_491 : entity work.gfmul
port map(
a=>a_4,
b=>"1001101011",
X=>mulr_4_491);

mulr_1_492<=a_1;
mulc_2_492 : entity work.gfmul
port map(
a=>a_2,
b=>"0011101010",
X=>mulr_2_492);

mulc_3_492 : entity work.gfmul
port map(
a=>a_3,
b=>"0011111001",
X=>mulr_3_492);

mulc_4_492 : entity work.gfmul
port map(
a=>a_4,
b=>"1101111100",
X=>mulr_4_492);

mulr_1_493<=a_1;
mulc_2_493 : entity work.gfmul
port map(
a=>a_2,
b=>"0111010100",
X=>mulr_2_493);

mulc_3_493 : entity work.gfmul
port map(
a=>a_3,
b=>"1111100100",
X=>mulr_3_493);

mulc_4_493 : entity work.gfmul
port map(
a=>a_4,
b=>"1111010110",
X=>mulr_4_493);

mulr_1_494<=a_1;
mulc_2_494 : entity work.gfmul
port map(
a=>a_2,
b=>"1110101000",
X=>mulr_2_494);

mulc_3_494 : entity work.gfmul
port map(
a=>a_3,
b=>"1110001011",
X=>mulr_3_494);

mulc_4_494 : entity work.gfmul
port map(
a=>a_4,
b=>"1010001111",
X=>mulr_4_494);

mulr_1_495<=a_1;
mulc_2_495 : entity work.gfmul
port map(
a=>a_2,
b=>"1101011001",
X=>mulr_2_495);

mulc_3_495 : entity work.gfmul
port map(
a=>a_3,
b=>"1000110111",
X=>mulr_3_495);

mulc_4_495 : entity work.gfmul
port map(
a=>a_4,
b=>"0001010101",
X=>mulr_4_495);

mulr_1_496<=a_1;
mulc_2_496 : entity work.gfmul
port map(
a=>a_2,
b=>"1010111011",
X=>mulr_2_496);

mulc_3_496 : entity work.gfmul
port map(
a=>a_3,
b=>"0011001110",
X=>mulr_3_496);

mulc_4_496 : entity work.gfmul
port map(
a=>a_4,
b=>"1010101000",
X=>mulr_4_496);

mulr_1_497<=a_1;
mulc_2_497 : entity work.gfmul
port map(
a=>a_2,
b=>"0101111111",
X=>mulr_2_497);

mulc_3_497 : entity work.gfmul
port map(
a=>a_3,
b=>"1100111000",
X=>mulr_3_497);

mulc_4_497 : entity work.gfmul
port map(
a=>a_4,
b=>"0101101101",
X=>mulr_4_497);

mulr_1_498<=a_1;
mulc_2_498 : entity work.gfmul
port map(
a=>a_2,
b=>"1011111110",
X=>mulr_2_498);

mulc_3_498 : entity work.gfmul
port map(
a=>a_3,
b=>"0011111011",
X=>mulr_3_498);

mulc_4_498 : entity work.gfmul
port map(
a=>a_4,
b=>"1101111010",
X=>mulr_4_498);

mulr_1_499<=a_1;
mulc_2_499 : entity work.gfmul
port map(
a=>a_2,
b=>"0111110101",
X=>mulr_2_499);

mulc_3_499 : entity work.gfmul
port map(
a=>a_3,
b=>"1111101100",
X=>mulr_3_499);

mulc_4_499 : entity work.gfmul
port map(
a=>a_4,
b=>"1111100110",
X=>mulr_4_499);

mulr_1_500<=a_1;
mulc_2_500 : entity work.gfmul
port map(
a=>a_2,
b=>"1111101010",
X=>mulr_2_500);

mulc_3_500 : entity work.gfmul
port map(
a=>a_3,
b=>"1110101011",
X=>mulr_3_500);

mulc_4_500 : entity work.gfmul
port map(
a=>a_4,
b=>"1100001111",
X=>mulr_4_500);

mulr_1_501<=a_1;
mulc_2_501 : entity work.gfmul
port map(
a=>a_2,
b=>"1111011101",
X=>mulr_2_501);

mulc_3_501 : entity work.gfmul
port map(
a=>a_3,
b=>"1010110111",
X=>mulr_3_501);

mulc_4_501 : entity work.gfmul
port map(
a=>a_4,
b=>"0001001110",
X=>mulr_4_501);

mulr_1_502<=a_1;
mulc_2_502 : entity work.gfmul
port map(
a=>a_2,
b=>"1110110011",
X=>mulr_2_502);

mulc_3_502 : entity work.gfmul
port map(
a=>a_3,
b=>"1011001110",
X=>mulr_3_502);

mulc_4_502 : entity work.gfmul
port map(
a=>a_4,
b=>"1001110000",
X=>mulr_4_502);

mulr_1_503<=a_1;
mulc_2_503 : entity work.gfmul
port map(
a=>a_2,
b=>"1101101111",
X=>mulr_2_503);

mulc_3_503 : entity work.gfmul
port map(
a=>a_3,
b=>"1100101010",
X=>mulr_3_503);

mulc_4_503 : entity work.gfmul
port map(
a=>a_4,
b=>"1110100100",
X=>mulr_4_503);

mulr_1_504<=a_1;
mulc_2_504 : entity work.gfmul
port map(
a=>a_2,
b=>"1011010111",
X=>mulr_2_504);

mulc_3_504 : entity work.gfmul
port map(
a=>a_3,
b=>"0010110011",
X=>mulr_3_504);

mulc_4_504 : entity work.gfmul
port map(
a=>a_4,
b=>"0100011111",
X=>mulr_4_504);

mulr_1_505<=a_1;
mulc_2_505 : entity work.gfmul
port map(
a=>a_2,
b=>"0110100111",
X=>mulr_2_505);

mulc_3_505 : entity work.gfmul
port map(
a=>a_3,
b=>"1011001100",
X=>mulr_3_505);

mulc_4_505 : entity work.gfmul
port map(
a=>a_4,
b=>"0011101010",
X=>mulr_4_505);

mulr_1_506<=a_1;
mulc_2_506 : entity work.gfmul
port map(
a=>a_2,
b=>"1101001110",
X=>mulr_2_506);

mulc_3_506 : entity work.gfmul
port map(
a=>a_3,
b=>"1100100010",
X=>mulr_3_506);

mulc_4_506 : entity work.gfmul
port map(
a=>a_4,
b=>"1101011001",
X=>mulr_4_506);

mulr_1_507<=a_1;
mulc_2_507 : entity work.gfmul
port map(
a=>a_2,
b=>"1010010101",
X=>mulr_2_507);

mulc_3_507 : entity work.gfmul
port map(
a=>a_3,
b=>"0010010011",
X=>mulr_3_507);

mulc_4_507 : entity work.gfmul
port map(
a=>a_4,
b=>"1011111110",
X=>mulr_4_507);

mulr_1_508<=a_1;
mulc_2_508 : entity work.gfmul
port map(
a=>a_2,
b=>"0100100011",
X=>mulr_2_508);

mulc_3_508 : entity work.gfmul
port map(
a=>a_3,
b=>"1001001100",
X=>mulr_3_508);

mulc_4_508 : entity work.gfmul
port map(
a=>a_4,
b=>"1111011101",
X=>mulr_4_508);

mulr_1_509<=a_1;
mulc_2_509 : entity work.gfmul
port map(
a=>a_2,
b=>"1001000110",
X=>mulr_2_509);

mulc_3_509 : entity work.gfmul
port map(
a=>a_3,
b=>"0100100010",
X=>mulr_3_509);

mulc_4_509 : entity work.gfmul
port map(
a=>a_4,
b=>"1011010111",
X=>mulr_4_509);

mulr_1_510<=a_1;
mulc_2_510 : entity work.gfmul
port map(
a=>a_2,
b=>"0010000101",
X=>mulr_2_510);

mulc_3_510 : entity work.gfmul
port map(
a=>a_3,
b=>"0010000001",
X=>mulr_3_510);

mulc_4_510 : entity work.gfmul
port map(
a=>a_4,
b=>"1010010101",
X=>mulr_4_510);

mulr_1_511<=a_1;
mulc_2_511 : entity work.gfmul
port map(
a=>a_2,
b=>"0100001010",
X=>mulr_2_511);

mulc_3_511 : entity work.gfmul
port map(
a=>a_3,
b=>"1000000100",
X=>mulr_3_511);

mulc_4_511 : entity work.gfmul
port map(
a=>a_4,
b=>"0010000101",
X=>mulr_4_511);

mulr_1_512<=a_1;
mulc_2_512 : entity work.gfmul
port map(
a=>a_2,
b=>"1000010100",
X=>mulr_2_512);

mulc_3_512 : entity work.gfmul
port map(
a=>a_3,
b=>"0000000010",
X=>mulr_3_512);

mulc_4_512 : entity work.gfmul
port map(
a=>a_4,
b=>"0000100001",
X=>mulr_4_512);

mulr_1_513<=a_1;
mulc_2_513 : entity work.gfmul
port map(
a=>a_2,
b=>"0000100001",
X=>mulr_2_513);

mulc_3_513 : entity work.gfmul
port map(
a=>a_3,
b=>"0000001000",
X=>mulr_3_513);

mulc_4_513 : entity work.gfmul
port map(
a=>a_4,
b=>"0100001000",
X=>mulr_4_513);

mulr_1_514<=a_1;
mulc_2_514 : entity work.gfmul
port map(
a=>a_2,
b=>"0001000010",
X=>mulr_2_514);

mulc_3_514 : entity work.gfmul
port map(
a=>a_3,
b=>"0000100000",
X=>mulr_3_514);

mulc_4_514 : entity work.gfmul
port map(
a=>a_4,
b=>"0001010010",
X=>mulr_4_514);

mulr_1_515<=a_1;
mulc_2_515 : entity work.gfmul
port map(
a=>a_2,
b=>"0010000100",
X=>mulr_2_515);

mulc_3_515 : entity work.gfmul
port map(
a=>a_3,
b=>"0010000000",
X=>mulr_3_515);

mulc_4_515 : entity work.gfmul
port map(
a=>a_4,
b=>"1010010000",
X=>mulr_4_515);

mulr_1_516<=a_1;
mulc_2_516 : entity work.gfmul
port map(
a=>a_2,
b=>"0100001000",
X=>mulr_2_516);

mulc_3_516 : entity work.gfmul
port map(
a=>a_3,
b=>"1000000000",
X=>mulr_3_516);

mulc_4_516 : entity work.gfmul
port map(
a=>a_4,
b=>"0010101101",
X=>mulr_4_516);

mulr_1_517<=a_1;
mulc_2_517 : entity work.gfmul
port map(
a=>a_2,
b=>"1000010000",
X=>mulr_2_517);

mulc_3_517 : entity work.gfmul
port map(
a=>a_3,
b=>"0000010010",
X=>mulr_3_517);

mulc_4_517 : entity work.gfmul
port map(
a=>a_4,
b=>"0101100001",
X=>mulr_4_517);

mulr_1_518<=a_1;
mulc_2_518 : entity work.gfmul
port map(
a=>a_2,
b=>"0000101001",
X=>mulr_2_518);

mulc_3_518 : entity work.gfmul
port map(
a=>a_3,
b=>"0001001000",
X=>mulr_3_518);

mulc_4_518 : entity work.gfmul
port map(
a=>a_4,
b=>"1100011010",
X=>mulr_4_518);

mulr_1_519<=a_1;
mulc_2_519 : entity work.gfmul
port map(
a=>a_2,
b=>"0001010010",
X=>mulr_2_519);

mulc_3_519 : entity work.gfmul
port map(
a=>a_3,
b=>"0100100000",
X=>mulr_3_519);

mulc_4_519 : entity work.gfmul
port map(
a=>a_4,
b=>"0011100110",
X=>mulr_4_519);

mulr_1_520<=a_1;
mulc_2_520 : entity work.gfmul
port map(
a=>a_2,
b=>"0010100100",
X=>mulr_2_520);

mulc_3_520 : entity work.gfmul
port map(
a=>a_3,
b=>"0010001001",
X=>mulr_3_520);

mulc_4_520 : entity work.gfmul
port map(
a=>a_4,
b=>"1100111001",
X=>mulr_4_520);

mulr_1_521<=a_1;
mulc_2_521 : entity work.gfmul
port map(
a=>a_2,
b=>"0101001000",
X=>mulr_2_521);

mulc_3_521 : entity work.gfmul
port map(
a=>a_3,
b=>"1000100100",
X=>mulr_3_521);

mulc_4_521 : entity work.gfmul
port map(
a=>a_4,
b=>"0111111110",
X=>mulr_4_521);

mulr_1_522<=a_1;
mulc_2_522 : entity work.gfmul
port map(
a=>a_2,
b=>"1010010000",
X=>mulr_2_522);

mulc_3_522 : entity work.gfmul
port map(
a=>a_3,
b=>"0010000010",
X=>mulr_3_522);

mulc_4_522 : entity work.gfmul
port map(
a=>a_4,
b=>"1111101011",
X=>mulr_4_522);

mulr_1_523<=a_1;
mulc_2_523 : entity work.gfmul
port map(
a=>a_2,
b=>"0100101001",
X=>mulr_2_523);

mulc_3_523 : entity work.gfmul
port map(
a=>a_3,
b=>"1000001000",
X=>mulr_3_523);

mulc_4_523 : entity work.gfmul
port map(
a=>a_4,
b=>"1101100111",
X=>mulr_4_523);

mulr_1_524<=a_1;
mulc_2_524 : entity work.gfmul
port map(
a=>a_2,
b=>"1001010010",
X=>mulr_2_524);

mulc_3_524 : entity work.gfmul
port map(
a=>a_3,
b=>"0000110010",
X=>mulr_3_524);

mulc_4_524 : entity work.gfmul
port map(
a=>a_4,
b=>"1100001110",
X=>mulr_4_524);

mulr_1_525<=a_1;
mulc_2_525 : entity work.gfmul
port map(
a=>a_2,
b=>"0010101101",
X=>mulr_2_525);

mulc_3_525 : entity work.gfmul
port map(
a=>a_3,
b=>"0011001000",
X=>mulr_3_525);

mulc_4_525 : entity work.gfmul
port map(
a=>a_4,
b=>"0001000110",
X=>mulr_4_525);

mulr_1_526<=a_1;
mulc_2_526 : entity work.gfmul
port map(
a=>a_2,
b=>"0101011010",
X=>mulr_2_526);

mulc_3_526 : entity work.gfmul
port map(
a=>a_3,
b=>"1100100000",
X=>mulr_3_526);

mulc_4_526 : entity work.gfmul
port map(
a=>a_4,
b=>"1000110000",
X=>mulr_4_526);

mulr_1_527<=a_1;
mulc_2_527 : entity work.gfmul
port map(
a=>a_2,
b=>"1010110100",
X=>mulr_2_527);

mulc_3_527 : entity work.gfmul
port map(
a=>a_3,
b=>"0010011011",
X=>mulr_3_527);

mulc_4_527 : entity work.gfmul
port map(
a=>a_4,
b=>"0110100100",
X=>mulr_4_527);

mulr_1_528<=a_1;
mulc_2_528 : entity work.gfmul
port map(
a=>a_2,
b=>"0101100001",
X=>mulr_2_528);

mulc_3_528 : entity work.gfmul
port map(
a=>a_3,
b=>"1001101100",
X=>mulr_3_528);

mulc_4_528 : entity work.gfmul
port map(
a=>a_4,
b=>"0100111011",
X=>mulr_4_528);

mulr_1_529<=a_1;
mulc_2_529 : entity work.gfmul
port map(
a=>a_2,
b=>"1011000010",
X=>mulr_2_529);

mulc_3_529 : entity work.gfmul
port map(
a=>a_3,
b=>"0110100010",
X=>mulr_3_529);

mulc_4_529 : entity work.gfmul
port map(
a=>a_4,
b=>"0111001010",
X=>mulr_4_529);

mulr_1_530<=a_1;
mulc_2_530 : entity work.gfmul
port map(
a=>a_2,
b=>"0110001101",
X=>mulr_2_530);

mulc_3_530 : entity work.gfmul
port map(
a=>a_3,
b=>"1010000001",
X=>mulr_3_530);

mulc_4_530 : entity work.gfmul
port map(
a=>a_4,
b=>"1001001011",
X=>mulr_4_530);

mulr_1_531<=a_1;
mulc_2_531 : entity work.gfmul
port map(
a=>a_2,
b=>"1100011010",
X=>mulr_2_531);

mulc_3_531 : entity work.gfmul
port map(
a=>a_3,
b=>"1000010110",
X=>mulr_3_531);

mulc_4_531 : entity work.gfmul
port map(
a=>a_4,
b=>"1001111100",
X=>mulr_4_531);

mulr_1_532<=a_1;
mulc_2_532 : entity work.gfmul
port map(
a=>a_2,
b=>"1000111101",
X=>mulr_2_532);

mulc_3_532 : entity work.gfmul
port map(
a=>a_3,
b=>"0001001010",
X=>mulr_3_532);

mulc_4_532 : entity work.gfmul
port map(
a=>a_4,
b=>"1111000100",
X=>mulr_4_532);

mulr_1_533<=a_1;
mulc_2_533 : entity work.gfmul
port map(
a=>a_2,
b=>"0001110011",
X=>mulr_2_533);

mulc_3_533 : entity work.gfmul
port map(
a=>a_3,
b=>"0100101000",
X=>mulr_3_533);

mulc_4_533 : entity work.gfmul
port map(
a=>a_4,
b=>"1000011111",
X=>mulr_4_533);

mulr_1_534<=a_1;
mulc_2_534 : entity work.gfmul
port map(
a=>a_2,
b=>"0011100110",
X=>mulr_2_534);

mulc_3_534 : entity work.gfmul
port map(
a=>a_3,
b=>"0010101001",
X=>mulr_3_534);

mulc_4_534 : entity work.gfmul
port map(
a=>a_4,
b=>"0011011100",
X=>mulr_4_534);

mulr_1_535<=a_1;
mulc_2_535 : entity work.gfmul
port map(
a=>a_2,
b=>"0111001100",
X=>mulr_2_535);

mulc_3_535 : entity work.gfmul
port map(
a=>a_3,
b=>"1010100100",
X=>mulr_3_535);

mulc_4_535 : entity work.gfmul
port map(
a=>a_4,
b=>"1011101001",
X=>mulr_4_535);

mulr_1_536<=a_1;
mulc_2_536 : entity work.gfmul
port map(
a=>a_2,
b=>"1110011000",
X=>mulr_2_536);

mulc_3_536 : entity work.gfmul
port map(
a=>a_3,
b=>"1010000010",
X=>mulr_3_536);

mulc_4_536 : entity work.gfmul
port map(
a=>a_4,
b=>"1101100101",
X=>mulr_4_536);

mulr_1_537<=a_1;
mulc_2_537 : entity work.gfmul
port map(
a=>a_2,
b=>"1100111001",
X=>mulr_2_537);

mulc_3_537 : entity work.gfmul
port map(
a=>a_3,
b=>"1000011010",
X=>mulr_3_537);

mulc_4_537 : entity work.gfmul
port map(
a=>a_4,
b=>"1100011110",
X=>mulr_4_537);

mulr_1_538<=a_1;
mulc_2_538 : entity work.gfmul
port map(
a=>a_2,
b=>"1001111011",
X=>mulr_2_538);

mulc_3_538 : entity work.gfmul
port map(
a=>a_3,
b=>"0001111010",
X=>mulr_3_538);

mulc_4_538 : entity work.gfmul
port map(
a=>a_4,
b=>"0011000110",
X=>mulr_4_538);

mulr_1_539<=a_1;
mulc_2_539 : entity work.gfmul
port map(
a=>a_2,
b=>"0011111111",
X=>mulr_2_539);

mulc_3_539 : entity work.gfmul
port map(
a=>a_3,
b=>"0111101000",
X=>mulr_3_539);

mulc_4_539 : entity work.gfmul
port map(
a=>a_4,
b=>"1000111001",
X=>mulr_4_539);

mulr_1_540<=a_1;
mulc_2_540 : entity work.gfmul
port map(
a=>a_2,
b=>"0111111110",
X=>mulr_2_540);

mulc_3_540 : entity work.gfmul
port map(
a=>a_3,
b=>"1110101001",
X=>mulr_3_540);

mulc_4_540 : entity work.gfmul
port map(
a=>a_4,
b=>"0111101100",
X=>mulr_4_540);

mulr_1_541<=a_1;
mulc_2_541 : entity work.gfmul
port map(
a=>a_2,
b=>"1111111100",
X=>mulr_2_541);

mulc_3_541 : entity work.gfmul
port map(
a=>a_3,
b=>"1010111111",
X=>mulr_3_541);

mulc_4_541 : entity work.gfmul
port map(
a=>a_4,
b=>"1101111011",
X=>mulr_4_541);

mulr_1_542<=a_1;
mulc_2_542 : entity work.gfmul
port map(
a=>a_2,
b=>"1111110001",
X=>mulr_2_542);

mulc_3_542 : entity work.gfmul
port map(
a=>a_3,
b=>"1011101110",
X=>mulr_3_542);

mulc_4_542 : entity work.gfmul
port map(
a=>a_4,
b=>"1111101110",
X=>mulr_4_542);

mulr_1_543<=a_1;
mulc_2_543 : entity work.gfmul
port map(
a=>a_2,
b=>"1111101011",
X=>mulr_2_543);

mulc_3_543 : entity work.gfmul
port map(
a=>a_3,
b=>"1110101010",
X=>mulr_3_543);

mulc_4_543 : entity work.gfmul
port map(
a=>a_4,
b=>"1101001111",
X=>mulr_4_543);

mulr_1_544<=a_1;
mulc_2_544 : entity work.gfmul
port map(
a=>a_2,
b=>"1111011111",
X=>mulr_2_544);

mulc_3_544 : entity work.gfmul
port map(
a=>a_3,
b=>"1010110011",
X=>mulr_3_544);

mulc_4_544 : entity work.gfmul
port map(
a=>a_4,
b=>"1001001110",
X=>mulr_4_544);

mulr_1_545<=a_1;
mulc_2_545 : entity work.gfmul
port map(
a=>a_2,
b=>"1110110111",
X=>mulr_2_545);

mulc_3_545 : entity work.gfmul
port map(
a=>a_3,
b=>"1011011110",
X=>mulr_3_545);

mulc_4_545 : entity work.gfmul
port map(
a=>a_4,
b=>"1001010100",
X=>mulr_4_545);

mulr_1_546<=a_1;
mulc_2_546 : entity work.gfmul
port map(
a=>a_2,
b=>"1101100111",
X=>mulr_2_546);

mulc_3_546 : entity work.gfmul
port map(
a=>a_3,
b=>"1101101010",
X=>mulr_3_546);

mulc_4_546 : entity work.gfmul
port map(
a=>a_4,
b=>"1010000100",
X=>mulr_4_546);

mulr_1_547<=a_1;
mulc_2_547 : entity work.gfmul
port map(
a=>a_2,
b=>"1011000111",
X=>mulr_2_547);

mulc_3_547 : entity work.gfmul
port map(
a=>a_3,
b=>"0110110011",
X=>mulr_3_547);

mulc_4_547 : entity work.gfmul
port map(
a=>a_4,
b=>"0000001101",
X=>mulr_4_547);

mulr_1_548<=a_1;
mulc_2_548 : entity work.gfmul
port map(
a=>a_2,
b=>"0110000111",
X=>mulr_2_548);

mulc_3_548 : entity work.gfmul
port map(
a=>a_3,
b=>"1011000101",
X=>mulr_3_548);

mulc_4_548 : entity work.gfmul
port map(
a=>a_4,
b=>"0001101000",
X=>mulr_4_548);

mulr_1_549<=a_1;
mulc_2_549 : entity work.gfmul
port map(
a=>a_2,
b=>"1100001110",
X=>mulr_2_549);

mulc_3_549 : entity work.gfmul
port map(
a=>a_3,
b=>"1100000110",
X=>mulr_3_549);

mulc_4_549 : entity work.gfmul
port map(
a=>a_4,
b=>"1101000000",
X=>mulr_4_549);

mulr_1_550<=a_1;
mulc_2_550 : entity work.gfmul
port map(
a=>a_2,
b=>"1000010101",
X=>mulr_2_550);

mulc_3_550 : entity work.gfmul
port map(
a=>a_3,
b=>"0000000011",
X=>mulr_3_550);

mulc_4_550 : entity work.gfmul
port map(
a=>a_4,
b=>"1000110110",
X=>mulr_4_550);

mulr_1_551<=a_1;
mulc_2_551 : entity work.gfmul
port map(
a=>a_2,
b=>"0000100011",
X=>mulr_2_551);

mulc_3_551 : entity work.gfmul
port map(
a=>a_3,
b=>"0000001100",
X=>mulr_3_551);

mulc_4_551 : entity work.gfmul
port map(
a=>a_4,
b=>"0110010100",
X=>mulr_4_551);

mulr_1_552<=a_1;
mulc_2_552 : entity work.gfmul
port map(
a=>a_2,
b=>"0001000110",
X=>mulr_2_552);

mulc_3_552 : entity work.gfmul
port map(
a=>a_3,
b=>"0000110000",
X=>mulr_3_552);

mulc_4_552 : entity work.gfmul
port map(
a=>a_4,
b=>"0010111011",
X=>mulr_4_552);

mulr_1_553<=a_1;
mulc_2_553 : entity work.gfmul
port map(
a=>a_2,
b=>"0010001100",
X=>mulr_2_553);

mulc_3_553 : entity work.gfmul
port map(
a=>a_3,
b=>"0011000000",
X=>mulr_3_553);

mulc_4_553 : entity work.gfmul
port map(
a=>a_4,
b=>"0111010001",
X=>mulr_4_553);

mulr_1_554<=a_1;
mulc_2_554 : entity work.gfmul
port map(
a=>a_2,
b=>"0100011000",
X=>mulr_2_554);

mulc_3_554 : entity work.gfmul
port map(
a=>a_3,
b=>"1100000000",
X=>mulr_3_554);

mulc_4_554 : entity work.gfmul
port map(
a=>a_4,
b=>"1010010011",
X=>mulr_4_554);

mulr_1_555<=a_1;
mulc_2_555 : entity work.gfmul
port map(
a=>a_2,
b=>"1000110000",
X=>mulr_2_555);

mulc_3_555 : entity work.gfmul
port map(
a=>a_3,
b=>"0000011011",
X=>mulr_3_555);

mulc_4_555 : entity work.gfmul
port map(
a=>a_4,
b=>"0010110101",
X=>mulr_4_555);

mulr_1_556<=a_1;
mulc_2_556 : entity work.gfmul
port map(
a=>a_2,
b=>"0001101001",
X=>mulr_2_556);

mulc_3_556 : entity work.gfmul
port map(
a=>a_3,
b=>"0001101100",
X=>mulr_3_556);

mulc_4_556 : entity work.gfmul
port map(
a=>a_4,
b=>"0110100001",
X=>mulr_4_556);

mulr_1_557<=a_1;
mulc_2_557 : entity work.gfmul
port map(
a=>a_2,
b=>"0011010010",
X=>mulr_2_557);

mulc_3_557 : entity work.gfmul
port map(
a=>a_3,
b=>"0110110000",
X=>mulr_3_557);

mulc_4_557 : entity work.gfmul
port map(
a=>a_4,
b=>"0100010011",
X=>mulr_4_557);

mulr_1_558<=a_1;
mulc_2_558 : entity work.gfmul
port map(
a=>a_2,
b=>"0110100100",
X=>mulr_2_558);

mulc_3_558 : entity work.gfmul
port map(
a=>a_3,
b=>"1011001001",
X=>mulr_3_558);

mulc_4_558 : entity work.gfmul
port map(
a=>a_4,
b=>"0010001010",
X=>mulr_4_558);

mulr_1_559<=a_1;
mulc_2_559 : entity work.gfmul
port map(
a=>a_2,
b=>"1101001000",
X=>mulr_2_559);

mulc_3_559 : entity work.gfmul
port map(
a=>a_3,
b=>"1100110110",
X=>mulr_3_559);

mulc_4_559 : entity work.gfmul
port map(
a=>a_4,
b=>"0001011001",
X=>mulr_4_559);

mulr_1_560<=a_1;
mulc_2_560 : entity work.gfmul
port map(
a=>a_2,
b=>"1010011001",
X=>mulr_2_560);

mulc_3_560 : entity work.gfmul
port map(
a=>a_3,
b=>"0011000011",
X=>mulr_3_560);

mulc_4_560 : entity work.gfmul
port map(
a=>a_4,
b=>"1011001000",
X=>mulr_4_560);

mulr_1_561<=a_1;
mulc_2_561 : entity work.gfmul
port map(
a=>a_2,
b=>"0100111011",
X=>mulr_2_561);

mulc_3_561 : entity work.gfmul
port map(
a=>a_3,
b=>"1100001100",
X=>mulr_3_561);

mulc_4_561 : entity work.gfmul
port map(
a=>a_4,
b=>"1001101101",
X=>mulr_4_561);

mulr_1_562<=a_1;
mulc_2_562 : entity work.gfmul
port map(
a=>a_2,
b=>"1001110110",
X=>mulr_2_562);

mulc_3_562 : entity work.gfmul
port map(
a=>a_3,
b=>"0000101011",
X=>mulr_3_562);

mulc_4_562 : entity work.gfmul
port map(
a=>a_4,
b=>"1101001100",
X=>mulr_4_562);

mulr_1_563<=a_1;
mulc_2_563 : entity work.gfmul
port map(
a=>a_2,
b=>"0011100101",
X=>mulr_2_563);

mulc_3_563 : entity work.gfmul
port map(
a=>a_3,
b=>"0010101100",
X=>mulr_3_563);

mulc_4_563 : entity work.gfmul
port map(
a=>a_4,
b=>"1001010110",
X=>mulr_4_563);

mulr_1_564<=a_1;
mulc_2_564 : entity work.gfmul
port map(
a=>a_2,
b=>"0111001010",
X=>mulr_2_564);

mulc_3_564 : entity work.gfmul
port map(
a=>a_3,
b=>"1010110000",
X=>mulr_3_564);

mulc_4_564 : entity work.gfmul
port map(
a=>a_4,
b=>"1010010100",
X=>mulr_4_564);

mulr_1_565<=a_1;
mulc_2_565 : entity work.gfmul
port map(
a=>a_2,
b=>"1110010100",
X=>mulr_2_565);

mulc_3_565 : entity work.gfmul
port map(
a=>a_3,
b=>"1011010010",
X=>mulr_3_565);

mulc_4_565 : entity work.gfmul
port map(
a=>a_4,
b=>"0010001101",
X=>mulr_4_565);

mulr_1_566<=a_1;
mulc_2_566 : entity work.gfmul
port map(
a=>a_2,
b=>"1100100001",
X=>mulr_2_566);

mulc_3_566 : entity work.gfmul
port map(
a=>a_3,
b=>"1101011010",
X=>mulr_3_566);

mulc_4_566 : entity work.gfmul
port map(
a=>a_4,
b=>"0001100001",
X=>mulr_4_566);

mulr_1_567<=a_1;
mulc_2_567 : entity work.gfmul
port map(
a=>a_2,
b=>"1001001011",
X=>mulr_2_567);

mulc_3_567 : entity work.gfmul
port map(
a=>a_3,
b=>"0101110011",
X=>mulr_3_567);

mulc_4_567 : entity work.gfmul
port map(
a=>a_4,
b=>"1100001000",
X=>mulr_4_567);

mulr_1_568<=a_1;
mulc_2_568 : entity work.gfmul
port map(
a=>a_2,
b=>"0010011111",
X=>mulr_2_568);

mulc_3_568 : entity work.gfmul
port map(
a=>a_3,
b=>"0111000101",
X=>mulr_3_568);

mulc_4_568 : entity work.gfmul
port map(
a=>a_4,
b=>"0001110110",
X=>mulr_4_568);

mulr_1_569<=a_1;
mulc_2_569 : entity work.gfmul
port map(
a=>a_2,
b=>"0100111110",
X=>mulr_2_569);

mulc_3_569 : entity work.gfmul
port map(
a=>a_3,
b=>"1100011101",
X=>mulr_3_569);

mulc_4_569 : entity work.gfmul
port map(
a=>a_4,
b=>"1110110000",
X=>mulr_4_569);

mulr_1_570<=a_1;
mulc_2_570 : entity work.gfmul
port map(
a=>a_2,
b=>"1001111100",
X=>mulr_2_570);

mulc_3_570 : entity work.gfmul
port map(
a=>a_3,
b=>"0001101111",
X=>mulr_3_570);

mulc_4_570 : entity work.gfmul
port map(
a=>a_4,
b=>"0110111111",
X=>mulr_4_570);

mulr_1_571<=a_1;
mulc_2_571 : entity work.gfmul
port map(
a=>a_2,
b=>"0011110001",
X=>mulr_2_571);

mulc_3_571 : entity work.gfmul
port map(
a=>a_3,
b=>"0110111100",
X=>mulr_3_571);

mulc_4_571 : entity work.gfmul
port map(
a=>a_4,
b=>"0111100011",
X=>mulr_4_571);

mulr_1_572<=a_1;
mulc_2_572 : entity work.gfmul
port map(
a=>a_2,
b=>"0111100010",
X=>mulr_2_572);

mulc_3_572 : entity work.gfmul
port map(
a=>a_3,
b=>"1011111001",
X=>mulr_3_572);

mulc_4_572 : entity work.gfmul
port map(
a=>a_4,
b=>"1100000011",
X=>mulr_4_572);

mulr_1_573<=a_1;
mulc_2_573 : entity work.gfmul
port map(
a=>a_2,
b=>"1111000100",
X=>mulr_2_573);

mulc_3_573 : entity work.gfmul
port map(
a=>a_3,
b=>"1111110110",
X=>mulr_3_573);

mulc_4_573 : entity work.gfmul
port map(
a=>a_4,
b=>"0000101110",
X=>mulr_4_573);

mulr_1_574<=a_1;
mulc_2_574 : entity work.gfmul
port map(
a=>a_2,
b=>"1110000001",
X=>mulr_2_574);

mulc_3_574 : entity work.gfmul
port map(
a=>a_3,
b=>"1111000011",
X=>mulr_3_574);

mulc_4_574 : entity work.gfmul
port map(
a=>a_4,
b=>"0101110000",
X=>mulr_4_574);

mulr_1_575<=a_1;
mulc_2_575 : entity work.gfmul
port map(
a=>a_2,
b=>"1100001011",
X=>mulr_2_575);

mulc_3_575 : entity work.gfmul
port map(
a=>a_3,
b=>"1100010111",
X=>mulr_3_575);

mulc_4_575 : entity work.gfmul
port map(
a=>a_4,
b=>"1110010010",
X=>mulr_4_575);

mulr_1_576<=a_1;
mulc_2_576 : entity work.gfmul
port map(
a=>a_2,
b=>"1000011111",
X=>mulr_2_576);

mulc_3_576 : entity work.gfmul
port map(
a=>a_3,
b=>"0001000111",
X=>mulr_3_576);

mulc_4_576 : entity work.gfmul
port map(
a=>a_4,
b=>"0010101111",
X=>mulr_4_576);

mulr_1_577<=a_1;
mulc_2_577 : entity work.gfmul
port map(
a=>a_2,
b=>"0000110111",
X=>mulr_2_577);

mulc_3_577 : entity work.gfmul
port map(
a=>a_3,
b=>"0100011100",
X=>mulr_3_577);

mulc_4_577 : entity work.gfmul
port map(
a=>a_4,
b=>"0101110001",
X=>mulr_4_577);

mulr_1_578<=a_1;
mulc_2_578 : entity work.gfmul
port map(
a=>a_2,
b=>"0001101110",
X=>mulr_2_578);

mulc_3_578 : entity work.gfmul
port map(
a=>a_3,
b=>"0001111001",
X=>mulr_3_578);

mulc_4_578 : entity work.gfmul
port map(
a=>a_4,
b=>"1110011010",
X=>mulr_4_578);

mulr_1_579<=a_1;
mulc_2_579 : entity work.gfmul
port map(
a=>a_2,
b=>"0011011100",
X=>mulr_2_579);

mulc_3_579 : entity work.gfmul
port map(
a=>a_3,
b=>"0111100100",
X=>mulr_3_579);

mulc_4_579 : entity work.gfmul
port map(
a=>a_4,
b=>"0011101111",
X=>mulr_4_579);

mulr_1_580<=a_1;
mulc_2_580 : entity work.gfmul
port map(
a=>a_2,
b=>"0110111000",
X=>mulr_2_580);

mulc_3_580 : entity work.gfmul
port map(
a=>a_3,
b=>"1110011001",
X=>mulr_3_580);

mulc_4_580 : entity work.gfmul
port map(
a=>a_4,
b=>"1101110001",
X=>mulr_4_580);

mulr_1_581<=a_1;
mulc_2_581 : entity work.gfmul
port map(
a=>a_2,
b=>"1101110000",
X=>mulr_2_581);

mulc_3_581 : entity work.gfmul
port map(
a=>a_3,
b=>"1001111111",
X=>mulr_3_581);

mulc_4_581 : entity work.gfmul
port map(
a=>a_4,
b=>"1110111110",
X=>mulr_4_581);

mulr_1_582<=a_1;
mulc_2_582 : entity work.gfmul
port map(
a=>a_2,
b=>"1011101001",
X=>mulr_2_582);

mulc_3_582 : entity work.gfmul
port map(
a=>a_3,
b=>"0111101110",
X=>mulr_3_582);

mulc_4_582 : entity work.gfmul
port map(
a=>a_4,
b=>"0111001111",
X=>mulr_4_582);

mulr_1_583<=a_1;
mulc_2_583 : entity work.gfmul
port map(
a=>a_2,
b=>"0111011011",
X=>mulr_2_583);

mulc_3_583 : entity work.gfmul
port map(
a=>a_3,
b=>"1110110001",
X=>mulr_3_583);

mulc_4_583 : entity work.gfmul
port map(
a=>a_4,
b=>"1001100011",
X=>mulr_4_583);

mulr_1_584<=a_1;
mulc_2_584 : entity work.gfmul
port map(
a=>a_2,
b=>"1110110110",
X=>mulr_2_584);

mulc_3_584 : entity work.gfmul
port map(
a=>a_3,
b=>"1011011111",
X=>mulr_3_584);

mulc_4_584 : entity work.gfmul
port map(
a=>a_4,
b=>"1100111100",
X=>mulr_4_584);

mulr_1_585<=a_1;
mulc_2_585 : entity work.gfmul
port map(
a=>a_2,
b=>"1101100101",
X=>mulr_2_585);

mulc_3_585 : entity work.gfmul
port map(
a=>a_3,
b=>"1101101110",
X=>mulr_3_585);

mulc_4_585 : entity work.gfmul
port map(
a=>a_4,
b=>"0111010110",
X=>mulr_4_585);

mulr_1_586<=a_1;
mulc_2_586 : entity work.gfmul
port map(
a=>a_2,
b=>"1011000011",
X=>mulr_2_586);

mulc_3_586 : entity work.gfmul
port map(
a=>a_3,
b=>"0110100011",
X=>mulr_3_586);

mulc_4_586 : entity work.gfmul
port map(
a=>a_4,
b=>"1010101011",
X=>mulr_4_586);

mulr_1_587<=a_1;
mulc_2_587 : entity work.gfmul
port map(
a=>a_2,
b=>"0110001111",
X=>mulr_2_587);

mulc_3_587 : entity work.gfmul
port map(
a=>a_3,
b=>"1010000101",
X=>mulr_3_587);

mulc_4_587 : entity work.gfmul
port map(
a=>a_4,
b=>"0101110101",
X=>mulr_4_587);

mulr_1_588<=a_1;
mulc_2_588 : entity work.gfmul
port map(
a=>a_2,
b=>"1100011110",
X=>mulr_2_588);

mulc_3_588 : entity work.gfmul
port map(
a=>a_3,
b=>"1000000110",
X=>mulr_3_588);

mulc_4_588 : entity work.gfmul
port map(
a=>a_4,
b=>"1110111010",
X=>mulr_4_588);

mulr_1_589<=a_1;
mulc_2_589 : entity work.gfmul
port map(
a=>a_2,
b=>"1000110101",
X=>mulr_2_589);

mulc_3_589 : entity work.gfmul
port map(
a=>a_3,
b=>"0000001010",
X=>mulr_3_589);

mulc_4_589 : entity work.gfmul
port map(
a=>a_4,
b=>"0111101111",
X=>mulr_4_589);

mulr_1_590<=a_1;
mulc_2_590 : entity work.gfmul
port map(
a=>a_2,
b=>"0001100011",
X=>mulr_2_590);

mulc_3_590 : entity work.gfmul
port map(
a=>a_3,
b=>"0000101000",
X=>mulr_3_590);

mulc_4_590 : entity work.gfmul
port map(
a=>a_4,
b=>"1101100011",
X=>mulr_4_590);

mulr_1_591<=a_1;
mulc_2_591 : entity work.gfmul
port map(
a=>a_2,
b=>"0011000110",
X=>mulr_2_591);

mulc_3_591 : entity work.gfmul
port map(
a=>a_3,
b=>"0010100000",
X=>mulr_3_591);

mulc_4_591 : entity work.gfmul
port map(
a=>a_4,
b=>"1100101110",
X=>mulr_4_591);

mulr_1_592<=a_1;
mulc_2_592 : entity work.gfmul
port map(
a=>a_2,
b=>"0110001100",
X=>mulr_2_592);

mulc_3_592 : entity work.gfmul
port map(
a=>a_3,
b=>"1010000000",
X=>mulr_3_592);

mulc_4_592 : entity work.gfmul
port map(
a=>a_4,
b=>"0101000110",
X=>mulr_4_592);

mulr_1_593<=a_1;
mulc_2_593 : entity work.gfmul
port map(
a=>a_2,
b=>"1100011000",
X=>mulr_2_593);

mulc_3_593 : entity work.gfmul
port map(
a=>a_3,
b=>"1000010010",
X=>mulr_3_593);

mulc_4_593 : entity work.gfmul
port map(
a=>a_4,
b=>"1000100010",
X=>mulr_4_593);

mulr_1_594<=a_1;
mulc_2_594 : entity work.gfmul
port map(
a=>a_2,
b=>"1000111001",
X=>mulr_2_594);

mulc_3_594 : entity work.gfmul
port map(
a=>a_3,
b=>"0001011010",
X=>mulr_3_594);

mulc_4_594 : entity work.gfmul
port map(
a=>a_4,
b=>"0100110100",
X=>mulr_4_594);

mulr_1_595<=a_1;
mulc_2_595 : entity work.gfmul
port map(
a=>a_2,
b=>"0001111011",
X=>mulr_2_595);

mulc_3_595 : entity work.gfmul
port map(
a=>a_3,
b=>"0101101000",
X=>mulr_3_595);

mulc_4_595 : entity work.gfmul
port map(
a=>a_4,
b=>"0110110010",
X=>mulr_4_595);

mulr_1_596<=a_1;
mulc_2_596 : entity work.gfmul
port map(
a=>a_2,
b=>"0011110110",
X=>mulr_2_596);

mulc_3_596 : entity work.gfmul
port map(
a=>a_3,
b=>"0110101001",
X=>mulr_3_596);

mulc_4_596 : entity work.gfmul
port map(
a=>a_4,
b=>"0110001011",
X=>mulr_4_596);

mulr_1_597<=a_1;
mulc_2_597 : entity work.gfmul
port map(
a=>a_2,
b=>"0111101100",
X=>mulr_2_597);

mulc_3_597 : entity work.gfmul
port map(
a=>a_3,
b=>"1010101101",
X=>mulr_3_597);

mulc_4_597 : entity work.gfmul
port map(
a=>a_4,
b=>"0001000011",
X=>mulr_4_597);

mulr_1_598<=a_1;
mulc_2_598 : entity work.gfmul
port map(
a=>a_2,
b=>"1111011000",
X=>mulr_2_598);

mulc_3_598 : entity work.gfmul
port map(
a=>a_3,
b=>"1010100110",
X=>mulr_3_598);

mulc_4_598 : entity work.gfmul
port map(
a=>a_4,
b=>"1000011000",
X=>mulr_4_598);

mulr_1_599<=a_1;
mulc_2_599 : entity work.gfmul
port map(
a=>a_2,
b=>"1110111001",
X=>mulr_2_599);

mulc_3_599 : entity work.gfmul
port map(
a=>a_3,
b=>"1010001010",
X=>mulr_3_599);

mulc_4_599 : entity work.gfmul
port map(
a=>a_4,
b=>"0011100100",
X=>mulr_4_599);

mulr_1_600<=a_1;
mulc_2_600 : entity work.gfmul
port map(
a=>a_2,
b=>"1101111011",
X=>mulr_2_600);

mulc_3_600 : entity work.gfmul
port map(
a=>a_3,
b=>"1000111010",
X=>mulr_3_600);

mulc_4_600 : entity work.gfmul
port map(
a=>a_4,
b=>"1100101001",
X=>mulr_4_600);

mulr_1_601<=a_1;
mulc_2_601 : entity work.gfmul
port map(
a=>a_2,
b=>"1011111111",
X=>mulr_2_601);

mulc_3_601 : entity work.gfmul
port map(
a=>a_3,
b=>"0011111010",
X=>mulr_3_601);

mulc_4_601 : entity work.gfmul
port map(
a=>a_4,
b=>"0101111110",
X=>mulr_4_601);

mulr_1_602<=a_1;
mulc_2_602 : entity work.gfmul
port map(
a=>a_2,
b=>"0111110111",
X=>mulr_2_602);

mulc_3_602 : entity work.gfmul
port map(
a=>a_3,
b=>"1111101000",
X=>mulr_3_602);

mulc_4_602 : entity work.gfmul
port map(
a=>a_4,
b=>"1111100010",
X=>mulr_4_602);

mulr_1_603<=a_1;
mulc_2_603 : entity work.gfmul
port map(
a=>a_2,
b=>"1111101110",
X=>mulr_2_603);

mulc_3_603 : entity work.gfmul
port map(
a=>a_3,
b=>"1110111011",
X=>mulr_3_603);

mulc_4_603 : entity work.gfmul
port map(
a=>a_4,
b=>"1100101111",
X=>mulr_4_603);

mulr_1_604<=a_1;
mulc_2_604 : entity work.gfmul
port map(
a=>a_2,
b=>"1111010101",
X=>mulr_2_604);

mulc_3_604 : entity work.gfmul
port map(
a=>a_3,
b=>"1011110111",
X=>mulr_3_604);

mulc_4_604 : entity work.gfmul
port map(
a=>a_4,
b=>"0101001110",
X=>mulr_4_604);

mulr_1_605<=a_1;
mulc_2_605 : entity work.gfmul
port map(
a=>a_2,
b=>"1110100011",
X=>mulr_2_605);

mulc_3_605 : entity work.gfmul
port map(
a=>a_3,
b=>"1111001110",
X=>mulr_3_605);

mulc_4_605 : entity work.gfmul
port map(
a=>a_4,
b=>"1001100010",
X=>mulr_4_605);

mulr_1_606<=a_1;
mulc_2_606 : entity work.gfmul
port map(
a=>a_2,
b=>"1101001111",
X=>mulr_2_606);

mulc_3_606 : entity work.gfmul
port map(
a=>a_3,
b=>"1100100011",
X=>mulr_3_606);

mulc_4_606 : entity work.gfmul
port map(
a=>a_4,
b=>"1100110100",
X=>mulr_4_606);

mulr_1_607<=a_1;
mulc_2_607 : entity work.gfmul
port map(
a=>a_2,
b=>"1010010111",
X=>mulr_2_607);

mulc_3_607 : entity work.gfmul
port map(
a=>a_3,
b=>"0010010111",
X=>mulr_3_607);

mulc_4_607 : entity work.gfmul
port map(
a=>a_4,
b=>"0110010110",
X=>mulr_4_607);

mulr_1_608<=a_1;
mulc_2_608 : entity work.gfmul
port map(
a=>a_2,
b=>"0100100111",
X=>mulr_2_608);

mulc_3_608 : entity work.gfmul
port map(
a=>a_3,
b=>"1001011100",
X=>mulr_3_608);

mulc_4_608 : entity work.gfmul
port map(
a=>a_4,
b=>"0010101011",
X=>mulr_4_608);

mulr_1_609<=a_1;
mulc_2_609 : entity work.gfmul
port map(
a=>a_2,
b=>"1001001110",
X=>mulr_2_609);

mulc_3_609 : entity work.gfmul
port map(
a=>a_3,
b=>"0101100010",
X=>mulr_3_609);

mulc_4_609 : entity work.gfmul
port map(
a=>a_4,
b=>"0101010001",
X=>mulr_4_609);

mulr_1_610<=a_1;
mulc_2_610 : entity work.gfmul
port map(
a=>a_2,
b=>"0010010101",
X=>mulr_2_610);

mulc_3_610 : entity work.gfmul
port map(
a=>a_3,
b=>"0110000001",
X=>mulr_3_610);

mulc_4_610 : entity work.gfmul
port map(
a=>a_4,
b=>"1010011010",
X=>mulr_4_610);

mulr_1_611<=a_1;
mulc_2_611 : entity work.gfmul
port map(
a=>a_2,
b=>"0100101010",
X=>mulr_2_611);

mulc_3_611 : entity work.gfmul
port map(
a=>a_3,
b=>"1000001101",
X=>mulr_3_611);

mulc_4_611 : entity work.gfmul
port map(
a=>a_4,
b=>"0011111101",
X=>mulr_4_611);

mulr_1_612<=a_1;
mulc_2_612 : entity work.gfmul
port map(
a=>a_2,
b=>"1001010100",
X=>mulr_2_612);

mulc_3_612 : entity work.gfmul
port map(
a=>a_3,
b=>"0000100110",
X=>mulr_3_612);

mulc_4_612 : entity work.gfmul
port map(
a=>a_4,
b=>"1111100001",
X=>mulr_4_612);

mulr_1_613<=a_1;
mulc_2_613 : entity work.gfmul
port map(
a=>a_2,
b=>"0010100001",
X=>mulr_2_613);

mulc_3_613 : entity work.gfmul
port map(
a=>a_3,
b=>"0010011000",
X=>mulr_3_613);

mulc_4_613 : entity work.gfmul
port map(
a=>a_4,
b=>"1100110111",
X=>mulr_4_613);

mulr_1_614<=a_1;
mulc_2_614 : entity work.gfmul
port map(
a=>a_2,
b=>"0101000010",
X=>mulr_2_614);

mulc_3_614 : entity work.gfmul
port map(
a=>a_3,
b=>"1001100000",
X=>mulr_3_614);

mulc_4_614 : entity work.gfmul
port map(
a=>a_4,
b=>"0110001110",
X=>mulr_4_614);

mulr_1_615<=a_1;
mulc_2_615 : entity work.gfmul
port map(
a=>a_2,
b=>"1010000100",
X=>mulr_2_615);

mulc_3_615 : entity work.gfmul
port map(
a=>a_3,
b=>"0110010010",
X=>mulr_3_615);

mulc_4_615 : entity work.gfmul
port map(
a=>a_4,
b=>"0001101011",
X=>mulr_4_615);

mulr_1_616<=a_1;
mulc_2_616 : entity work.gfmul
port map(
a=>a_2,
b=>"0100000001",
X=>mulr_2_616);

mulc_3_616 : entity work.gfmul
port map(
a=>a_3,
b=>"1001000001",
X=>mulr_3_616);

mulc_4_616 : entity work.gfmul
port map(
a=>a_4,
b=>"1101011000",
X=>mulr_4_616);

mulr_1_617<=a_1;
mulc_2_617 : entity work.gfmul
port map(
a=>a_2,
b=>"1000000010",
X=>mulr_2_617);

mulc_3_617 : entity work.gfmul
port map(
a=>a_3,
b=>"0100010110",
X=>mulr_3_617);

mulc_4_617 : entity work.gfmul
port map(
a=>a_4,
b=>"1011110110",
X=>mulr_4_617);

mulr_1_618<=a_1;
mulc_2_618 : entity work.gfmul
port map(
a=>a_2,
b=>"0000001101",
X=>mulr_2_618);

mulc_3_618 : entity work.gfmul
port map(
a=>a_3,
b=>"0001010001",
X=>mulr_3_618);

mulc_4_618 : entity work.gfmul
port map(
a=>a_4,
b=>"1110011101",
X=>mulr_4_618);

mulr_1_619<=a_1;
mulc_2_619 : entity work.gfmul
port map(
a=>a_2,
b=>"0000011010",
X=>mulr_2_619);

mulc_3_619 : entity work.gfmul
port map(
a=>a_3,
b=>"0101000100",
X=>mulr_3_619);

mulc_4_619 : entity work.gfmul
port map(
a=>a_4,
b=>"0011010111",
X=>mulr_4_619);

mulr_1_620<=a_1;
mulc_2_620 : entity work.gfmul
port map(
a=>a_2,
b=>"0000110100",
X=>mulr_2_620);

mulc_3_620 : entity work.gfmul
port map(
a=>a_3,
b=>"0100011001",
X=>mulr_3_620);

mulc_4_620 : entity work.gfmul
port map(
a=>a_4,
b=>"1010110001",
X=>mulr_4_620);

mulr_1_621<=a_1;
mulc_2_621 : entity work.gfmul
port map(
a=>a_2,
b=>"0001101000",
X=>mulr_2_621);

mulc_3_621 : entity work.gfmul
port map(
a=>a_3,
b=>"0001101101",
X=>mulr_3_621);

mulc_4_621 : entity work.gfmul
port map(
a=>a_4,
b=>"0110100101",
X=>mulr_4_621);

mulr_1_622<=a_1;
mulc_2_622 : entity work.gfmul
port map(
a=>a_2,
b=>"0011010000",
X=>mulr_2_622);

mulc_3_622 : entity work.gfmul
port map(
a=>a_3,
b=>"0110110100",
X=>mulr_3_622);

mulc_4_622 : entity work.gfmul
port map(
a=>a_4,
b=>"0100110011",
X=>mulr_4_622);

mulr_1_623<=a_1;
mulc_2_623 : entity work.gfmul
port map(
a=>a_2,
b=>"0110100000",
X=>mulr_2_623);

mulc_3_623 : entity work.gfmul
port map(
a=>a_3,
b=>"1011011001",
X=>mulr_3_623);

mulc_4_623 : entity work.gfmul
port map(
a=>a_4,
b=>"0110001010",
X=>mulr_4_623);

mulr_1_624<=a_1;
mulc_2_624 : entity work.gfmul
port map(
a=>a_2,
b=>"1101000000",
X=>mulr_2_624);

mulc_3_624 : entity work.gfmul
port map(
a=>a_3,
b=>"1101110110",
X=>mulr_3_624);

mulc_4_624 : entity work.gfmul
port map(
a=>a_4,
b=>"0001001011",
X=>mulr_4_624);

mulr_1_625<=a_1;
mulc_2_625 : entity work.gfmul
port map(
a=>a_2,
b=>"1010001001",
X=>mulr_2_625);

mulc_3_625 : entity work.gfmul
port map(
a=>a_3,
b=>"0111000011",
X=>mulr_3_625);

mulc_4_625 : entity work.gfmul
port map(
a=>a_4,
b=>"1001011000",
X=>mulr_4_625);

mulr_1_626<=a_1;
mulc_2_626 : entity work.gfmul
port map(
a=>a_2,
b=>"0100011011",
X=>mulr_2_626);

mulc_3_626 : entity work.gfmul
port map(
a=>a_3,
b=>"1100000101",
X=>mulr_3_626);

mulc_4_626 : entity work.gfmul
port map(
a=>a_4,
b=>"1011100100",
X=>mulr_4_626);

mulr_1_627<=a_1;
mulc_2_627 : entity work.gfmul
port map(
a=>a_2,
b=>"1000110110",
X=>mulr_2_627);

mulc_3_627 : entity work.gfmul
port map(
a=>a_3,
b=>"0000001111",
X=>mulr_3_627);

mulc_4_627 : entity work.gfmul
port map(
a=>a_4,
b=>"1100001101",
X=>mulr_4_627);

mulr_1_628<=a_1;
mulc_2_628 : entity work.gfmul
port map(
a=>a_2,
b=>"0001100101",
X=>mulr_2_628);

mulc_3_628 : entity work.gfmul
port map(
a=>a_3,
b=>"0000111100",
X=>mulr_3_628);

mulc_4_628 : entity work.gfmul
port map(
a=>a_4,
b=>"0001011110",
X=>mulr_4_628);

mulr_1_629<=a_1;
mulc_2_629 : entity work.gfmul
port map(
a=>a_2,
b=>"0011001010",
X=>mulr_2_629);

mulc_3_629 : entity work.gfmul
port map(
a=>a_3,
b=>"0011110000",
X=>mulr_3_629);

mulc_4_629 : entity work.gfmul
port map(
a=>a_4,
b=>"1011110000",
X=>mulr_4_629);

mulr_1_630<=a_1;
mulc_2_630 : entity work.gfmul
port map(
a=>a_2,
b=>"0110010100",
X=>mulr_2_630);

mulc_3_630 : entity work.gfmul
port map(
a=>a_3,
b=>"1111000000",
X=>mulr_3_630);

mulc_4_630 : entity work.gfmul
port map(
a=>a_4,
b=>"1110101101",
X=>mulr_4_630);

mulr_1_631<=a_1;
mulc_2_631 : entity work.gfmul
port map(
a=>a_2,
b=>"1100101000",
X=>mulr_2_631);

mulc_3_631 : entity work.gfmul
port map(
a=>a_3,
b=>"1100011011",
X=>mulr_3_631);

mulc_4_631 : entity work.gfmul
port map(
a=>a_4,
b=>"0101010111",
X=>mulr_4_631);

mulr_1_632<=a_1;
mulc_2_632 : entity work.gfmul
port map(
a=>a_2,
b=>"1001011001",
X=>mulr_2_632);

mulc_3_632 : entity work.gfmul
port map(
a=>a_3,
b=>"0001110111",
X=>mulr_3_632);

mulc_4_632 : entity work.gfmul
port map(
a=>a_4,
b=>"1010101010",
X=>mulr_4_632);

mulr_1_633<=a_1;
mulc_2_633 : entity work.gfmul
port map(
a=>a_2,
b=>"0010111011",
X=>mulr_2_633);

mulc_3_633 : entity work.gfmul
port map(
a=>a_3,
b=>"0111011100",
X=>mulr_3_633);

mulc_4_633 : entity work.gfmul
port map(
a=>a_4,
b=>"0101111101",
X=>mulr_4_633);

mulr_1_634<=a_1;
mulc_2_634 : entity work.gfmul
port map(
a=>a_2,
b=>"0101110110",
X=>mulr_2_634);

mulc_3_634 : entity work.gfmul
port map(
a=>a_3,
b=>"1101111001",
X=>mulr_3_634);

mulc_4_634 : entity work.gfmul
port map(
a=>a_4,
b=>"1111111010",
X=>mulr_4_634);

mulr_1_635<=a_1;
mulc_2_635 : entity work.gfmul
port map(
a=>a_2,
b=>"1011101100",
X=>mulr_2_635);

mulc_3_635 : entity work.gfmul
port map(
a=>a_3,
b=>"0111111111",
X=>mulr_3_635);

mulc_4_635 : entity work.gfmul
port map(
a=>a_4,
b=>"1111101111",
X=>mulr_4_635);

mulr_1_636<=a_1;
mulc_2_636 : entity work.gfmul
port map(
a=>a_2,
b=>"0111010001",
X=>mulr_2_636);

mulc_3_636 : entity work.gfmul
port map(
a=>a_3,
b=>"1111110101",
X=>mulr_3_636);

mulc_4_636 : entity work.gfmul
port map(
a=>a_4,
b=>"1101000111",
X=>mulr_4_636);

mulr_1_637<=a_1;
mulc_2_637 : entity work.gfmul
port map(
a=>a_2,
b=>"1110100010",
X=>mulr_2_637);

mulc_3_637 : entity work.gfmul
port map(
a=>a_3,
b=>"1111001111",
X=>mulr_3_637);

mulc_4_637 : entity work.gfmul
port map(
a=>a_4,
b=>"1000001110",
X=>mulr_4_637);

mulr_1_638<=a_1;
mulc_2_638 : entity work.gfmul
port map(
a=>a_2,
b=>"1101001101",
X=>mulr_2_638);

mulc_3_638 : entity work.gfmul
port map(
a=>a_3,
b=>"1100100111",
X=>mulr_3_638);

mulc_4_638 : entity work.gfmul
port map(
a=>a_4,
b=>"0001010100",
X=>mulr_4_638);

mulr_1_639<=a_1;
mulc_2_639 : entity work.gfmul
port map(
a=>a_2,
b=>"1010010011",
X=>mulr_2_639);

mulc_3_639 : entity work.gfmul
port map(
a=>a_3,
b=>"0010000111",
X=>mulr_3_639);

mulc_4_639 : entity work.gfmul
port map(
a=>a_4,
b=>"1010100000",
X=>mulr_4_639);

mulr_1_640<=a_1;
mulc_2_640 : entity work.gfmul
port map(
a=>a_2,
b=>"0100101111",
X=>mulr_2_640);

mulc_3_640 : entity work.gfmul
port map(
a=>a_3,
b=>"1000011100",
X=>mulr_3_640);

mulc_4_640 : entity work.gfmul
port map(
a=>a_4,
b=>"0100101101",
X=>mulr_4_640);

mulr_1_641<=a_1;
mulc_2_641 : entity work.gfmul
port map(
a=>a_2,
b=>"1001011110",
X=>mulr_2_641);

mulc_3_641 : entity work.gfmul
port map(
a=>a_3,
b=>"0001100010",
X=>mulr_3_641);

mulc_4_641 : entity work.gfmul
port map(
a=>a_4,
b=>"0101111010",
X=>mulr_4_641);

mulr_1_642<=a_1;
mulc_2_642 : entity work.gfmul
port map(
a=>a_2,
b=>"0010110101",
X=>mulr_2_642);

mulc_3_642 : entity work.gfmul
port map(
a=>a_3,
b=>"0110001000",
X=>mulr_3_642);

mulc_4_642 : entity work.gfmul
port map(
a=>a_4,
b=>"1111000010",
X=>mulr_4_642);

mulr_1_643<=a_1;
mulc_2_643 : entity work.gfmul
port map(
a=>a_2,
b=>"0101101010",
X=>mulr_2_643);

mulc_3_643 : entity work.gfmul
port map(
a=>a_3,
b=>"1000101001",
X=>mulr_3_643);

mulc_4_643 : entity work.gfmul
port map(
a=>a_4,
b=>"1000101111",
X=>mulr_4_643);

mulr_1_644<=a_1;
mulc_2_644 : entity work.gfmul
port map(
a=>a_2,
b=>"1011010100",
X=>mulr_2_644);

mulc_3_644 : entity work.gfmul
port map(
a=>a_3,
b=>"0010110110",
X=>mulr_3_644);

mulc_4_644 : entity work.gfmul
port map(
a=>a_4,
b=>"0101011100",
X=>mulr_4_644);

mulr_1_645<=a_1;
mulc_2_645 : entity work.gfmul
port map(
a=>a_2,
b=>"0110100001",
X=>mulr_2_645);

mulc_3_645 : entity work.gfmul
port map(
a=>a_3,
b=>"1011011000",
X=>mulr_3_645);

mulc_4_645 : entity work.gfmul
port map(
a=>a_4,
b=>"1011110010",
X=>mulr_4_645);

mulr_1_646<=a_1;
mulc_2_646 : entity work.gfmul
port map(
a=>a_2,
b=>"1101000010",
X=>mulr_2_646);

mulc_3_646 : entity work.gfmul
port map(
a=>a_3,
b=>"1101110010",
X=>mulr_3_646);

mulc_4_646 : entity work.gfmul
port map(
a=>a_4,
b=>"1110111101",
X=>mulr_4_646);

mulr_1_647<=a_1;
mulc_2_647 : entity work.gfmul
port map(
a=>a_2,
b=>"1010001101",
X=>mulr_2_647);

mulc_3_647 : entity work.gfmul
port map(
a=>a_3,
b=>"0111010011",
X=>mulr_3_647);

mulc_4_647 : entity work.gfmul
port map(
a=>a_4,
b=>"0111010111",
X=>mulr_4_647);

mulr_1_648<=a_1;
mulc_2_648 : entity work.gfmul
port map(
a=>a_2,
b=>"0100010011",
X=>mulr_2_648);

mulc_3_648 : entity work.gfmul
port map(
a=>a_3,
b=>"1101000101",
X=>mulr_3_648);

mulc_4_648 : entity work.gfmul
port map(
a=>a_4,
b=>"1010100011",
X=>mulr_4_648);

mulr_1_649<=a_1;
mulc_2_649 : entity work.gfmul
port map(
a=>a_2,
b=>"1000100110",
X=>mulr_2_649);

mulc_3_649 : entity work.gfmul
port map(
a=>a_3,
b=>"0100001111",
X=>mulr_3_649);

mulc_4_649 : entity work.gfmul
port map(
a=>a_4,
b=>"0100110101",
X=>mulr_4_649);

mulr_1_650<=a_1;
mulc_2_650 : entity work.gfmul
port map(
a=>a_2,
b=>"0001000101",
X=>mulr_2_650);

mulc_3_650 : entity work.gfmul
port map(
a=>a_3,
b=>"0000110101",
X=>mulr_3_650);

mulc_4_650 : entity work.gfmul
port map(
a=>a_4,
b=>"0110111010",
X=>mulr_4_650);

mulr_1_651<=a_1;
mulc_2_651 : entity work.gfmul
port map(
a=>a_2,
b=>"0010001010",
X=>mulr_2_651);

mulc_3_651 : entity work.gfmul
port map(
a=>a_3,
b=>"0011010100",
X=>mulr_3_651);

mulc_4_651 : entity work.gfmul
port map(
a=>a_4,
b=>"0111001011",
X=>mulr_4_651);

mulr_1_652<=a_1;
mulc_2_652 : entity work.gfmul
port map(
a=>a_2,
b=>"0100010100",
X=>mulr_2_652);

mulc_3_652 : entity work.gfmul
port map(
a=>a_3,
b=>"1101010000",
X=>mulr_3_652);

mulc_4_652 : entity work.gfmul
port map(
a=>a_4,
b=>"1001000011",
X=>mulr_4_652);

mulr_1_653<=a_1;
mulc_2_653 : entity work.gfmul
port map(
a=>a_2,
b=>"1000101000",
X=>mulr_2_653);

mulc_3_653 : entity work.gfmul
port map(
a=>a_3,
b=>"0101011011",
X=>mulr_3_653);

mulc_4_653 : entity work.gfmul
port map(
a=>a_4,
b=>"1000111100",
X=>mulr_4_653);

mulr_1_654<=a_1;
mulc_2_654 : entity work.gfmul
port map(
a=>a_2,
b=>"0001011001",
X=>mulr_2_654);

mulc_3_654 : entity work.gfmul
port map(
a=>a_3,
b=>"0101100101",
X=>mulr_3_654);

mulc_4_654 : entity work.gfmul
port map(
a=>a_4,
b=>"0111000100",
X=>mulr_4_654);

mulr_1_655<=a_1;
mulc_2_655 : entity work.gfmul
port map(
a=>a_2,
b=>"0010110010",
X=>mulr_2_655);

mulc_3_655 : entity work.gfmul
port map(
a=>a_3,
b=>"0110011101",
X=>mulr_3_655);

mulc_4_655 : entity work.gfmul
port map(
a=>a_4,
b=>"1000111011",
X=>mulr_4_655);

mulr_1_656<=a_1;
mulc_2_656 : entity work.gfmul
port map(
a=>a_2,
b=>"0101100100",
X=>mulr_2_656);

mulc_3_656 : entity work.gfmul
port map(
a=>a_3,
b=>"1001111101",
X=>mulr_3_656);

mulc_4_656 : entity work.gfmul
port map(
a=>a_4,
b=>"0111111100",
X=>mulr_4_656);

mulr_1_657<=a_1;
mulc_2_657 : entity work.gfmul
port map(
a=>a_2,
b=>"1011001000",
X=>mulr_2_657);

mulc_3_657 : entity work.gfmul
port map(
a=>a_3,
b=>"0111100110",
X=>mulr_3_657);

mulc_4_657 : entity work.gfmul
port map(
a=>a_4,
b=>"1111111011",
X=>mulr_4_657);

mulr_1_658<=a_1;
mulc_2_658 : entity work.gfmul
port map(
a=>a_2,
b=>"0110011001",
X=>mulr_2_658);

mulc_3_658 : entity work.gfmul
port map(
a=>a_3,
b=>"1110010001",
X=>mulr_3_658);

mulc_4_658 : entity work.gfmul
port map(
a=>a_4,
b=>"1111100111",
X=>mulr_4_658);

mulr_1_659<=a_1;
mulc_2_659 : entity work.gfmul
port map(
a=>a_2,
b=>"1100110010",
X=>mulr_2_659);

mulc_3_659 : entity work.gfmul
port map(
a=>a_3,
b=>"1001011111",
X=>mulr_3_659);

mulc_4_659 : entity work.gfmul
port map(
a=>a_4,
b=>"1100000111",
X=>mulr_4_659);

mulr_1_660<=a_1;
mulc_2_660 : entity work.gfmul
port map(
a=>a_2,
b=>"1001101101",
X=>mulr_2_660);

mulc_3_660 : entity work.gfmul
port map(
a=>a_3,
b=>"0101101110",
X=>mulr_3_660);

mulc_4_660 : entity work.gfmul
port map(
a=>a_4,
b=>"0000001110",
X=>mulr_4_660);

mulr_1_661<=a_1;
mulc_2_661 : entity work.gfmul
port map(
a=>a_2,
b=>"0011010011",
X=>mulr_2_661);

mulc_3_661 : entity work.gfmul
port map(
a=>a_3,
b=>"0110110001",
X=>mulr_3_661);

mulc_4_661 : entity work.gfmul
port map(
a=>a_4,
b=>"0001110000",
X=>mulr_4_661);

mulr_1_662<=a_1;
mulc_2_662 : entity work.gfmul
port map(
a=>a_2,
b=>"0110100110",
X=>mulr_2_662);

mulc_3_662 : entity work.gfmul
port map(
a=>a_3,
b=>"1011001101",
X=>mulr_3_662);

mulc_4_662 : entity work.gfmul
port map(
a=>a_4,
b=>"1110000000",
X=>mulr_4_662);

mulr_1_663<=a_1;
mulc_2_663 : entity work.gfmul
port map(
a=>a_2,
b=>"1101001100",
X=>mulr_2_663);

mulc_3_663 : entity work.gfmul
port map(
a=>a_3,
b=>"1100100110",
X=>mulr_3_663);

mulc_4_663 : entity work.gfmul
port map(
a=>a_4,
b=>"0000111111",
X=>mulr_4_663);

mulr_1_664<=a_1;
mulc_2_664 : entity work.gfmul
port map(
a=>a_2,
b=>"1010010001",
X=>mulr_2_664);

mulc_3_664 : entity work.gfmul
port map(
a=>a_3,
b=>"0010000011",
X=>mulr_3_664);

mulc_4_664 : entity work.gfmul
port map(
a=>a_4,
b=>"0111111000",
X=>mulr_4_664);

mulr_1_665<=a_1;
mulc_2_665 : entity work.gfmul
port map(
a=>a_2,
b=>"0100101011",
X=>mulr_2_665);

mulc_3_665 : entity work.gfmul
port map(
a=>a_3,
b=>"1000001100",
X=>mulr_3_665);

mulc_4_665 : entity work.gfmul
port map(
a=>a_4,
b=>"1111011011",
X=>mulr_4_665);

mulr_1_666<=a_1;
mulc_2_666 : entity work.gfmul
port map(
a=>a_2,
b=>"1001010110",
X=>mulr_2_666);

mulc_3_666 : entity work.gfmul
port map(
a=>a_3,
b=>"0000100010",
X=>mulr_3_666);

mulc_4_666 : entity work.gfmul
port map(
a=>a_4,
b=>"1011100111",
X=>mulr_4_666);

mulr_1_667<=a_1;
mulc_2_667 : entity work.gfmul
port map(
a=>a_2,
b=>"0010100101",
X=>mulr_2_667);

mulc_3_667 : entity work.gfmul
port map(
a=>a_3,
b=>"0010001000",
X=>mulr_3_667);

mulc_4_667 : entity work.gfmul
port map(
a=>a_4,
b=>"1100010101",
X=>mulr_4_667);

mulr_1_668<=a_1;
mulc_2_668 : entity work.gfmul
port map(
a=>a_2,
b=>"0101001010",
X=>mulr_2_668);

mulc_3_668 : entity work.gfmul
port map(
a=>a_3,
b=>"1000100000",
X=>mulr_3_668);

mulc_4_668 : entity work.gfmul
port map(
a=>a_4,
b=>"0010011110",
X=>mulr_4_668);

mulr_1_669<=a_1;
mulc_2_669 : entity work.gfmul
port map(
a=>a_2,
b=>"1010010100",
X=>mulr_2_669);

mulc_3_669 : entity work.gfmul
port map(
a=>a_3,
b=>"0010010010",
X=>mulr_3_669);

mulc_4_669 : entity work.gfmul
port map(
a=>a_4,
b=>"0011111001",
X=>mulr_4_669);

mulr_1_670<=a_1;
mulc_2_670 : entity work.gfmul
port map(
a=>a_2,
b=>"0100100001",
X=>mulr_2_670);

mulc_3_670 : entity work.gfmul
port map(
a=>a_3,
b=>"1001001000",
X=>mulr_3_670);

mulc_4_670 : entity work.gfmul
port map(
a=>a_4,
b=>"1111000001",
X=>mulr_4_670);

mulr_1_671<=a_1;
mulc_2_671 : entity work.gfmul
port map(
a=>a_2,
b=>"1001000010",
X=>mulr_2_671);

mulc_3_671 : entity work.gfmul
port map(
a=>a_3,
b=>"0100110010",
X=>mulr_3_671);

mulc_4_671 : entity work.gfmul
port map(
a=>a_4,
b=>"1000110111",
X=>mulr_4_671);

mulr_1_672<=a_1;
mulc_2_672 : entity work.gfmul
port map(
a=>a_2,
b=>"0010001101",
X=>mulr_2_672);

mulc_3_672 : entity work.gfmul
port map(
a=>a_3,
b=>"0011000001",
X=>mulr_3_672);

mulc_4_672 : entity work.gfmul
port map(
a=>a_4,
b=>"0110011100",
X=>mulr_4_672);

mulr_1_673<=a_1;
mulc_2_673 : entity work.gfmul
port map(
a=>a_2,
b=>"0100011010",
X=>mulr_2_673);

mulc_3_673 : entity work.gfmul
port map(
a=>a_3,
b=>"1100000100",
X=>mulr_3_673);

mulc_4_673 : entity work.gfmul
port map(
a=>a_4,
b=>"0011111011",
X=>mulr_4_673);

mulr_1_674<=a_1;
mulc_2_674 : entity work.gfmul
port map(
a=>a_2,
b=>"1000110100",
X=>mulr_2_674);

mulc_3_674 : entity work.gfmul
port map(
a=>a_3,
b=>"0000001011",
X=>mulr_3_674);

mulc_4_674 : entity work.gfmul
port map(
a=>a_4,
b=>"1111010001",
X=>mulr_4_674);

mulr_1_675<=a_1;
mulc_2_675 : entity work.gfmul
port map(
a=>a_2,
b=>"0001100001",
X=>mulr_2_675);

mulc_3_675 : entity work.gfmul
port map(
a=>a_3,
b=>"0000101100",
X=>mulr_3_675);

mulc_4_675 : entity work.gfmul
port map(
a=>a_4,
b=>"1010110111",
X=>mulr_4_675);

mulr_1_676<=a_1;
mulc_2_676 : entity work.gfmul
port map(
a=>a_2,
b=>"0011000010",
X=>mulr_2_676);

mulc_3_676 : entity work.gfmul
port map(
a=>a_3,
b=>"0010110000",
X=>mulr_3_676);

mulc_4_676 : entity work.gfmul
port map(
a=>a_4,
b=>"0110010101",
X=>mulr_4_676);

mulr_1_677<=a_1;
mulc_2_677 : entity work.gfmul
port map(
a=>a_2,
b=>"0110000100",
X=>mulr_2_677);

mulc_3_677 : entity work.gfmul
port map(
a=>a_3,
b=>"1011000000",
X=>mulr_3_677);

mulc_4_677 : entity work.gfmul
port map(
a=>a_4,
b=>"0010110011",
X=>mulr_4_677);

mulr_1_678<=a_1;
mulc_2_678 : entity work.gfmul
port map(
a=>a_2,
b=>"1100001000",
X=>mulr_2_678);

mulc_3_678 : entity work.gfmul
port map(
a=>a_3,
b=>"1100010010",
X=>mulr_3_678);

mulc_4_678 : entity work.gfmul
port map(
a=>a_4,
b=>"0110010001",
X=>mulr_4_678);

mulr_1_679<=a_1;
mulc_2_679 : entity work.gfmul
port map(
a=>a_2,
b=>"1000011001",
X=>mulr_2_679);

mulc_3_679 : entity work.gfmul
port map(
a=>a_3,
b=>"0001010011",
X=>mulr_3_679);

mulc_4_679 : entity work.gfmul
port map(
a=>a_4,
b=>"0010010011",
X=>mulr_4_679);

mulr_1_680<=a_1;
mulc_2_680 : entity work.gfmul
port map(
a=>a_2,
b=>"0000111011",
X=>mulr_2_680);

mulc_3_680 : entity work.gfmul
port map(
a=>a_3,
b=>"0101001100",
X=>mulr_3_680);

mulc_4_680 : entity work.gfmul
port map(
a=>a_4,
b=>"0010010001",
X=>mulr_4_680);

mulr_1_681<=a_1;
mulc_2_681 : entity work.gfmul
port map(
a=>a_2,
b=>"0001110110",
X=>mulr_2_681);

mulc_3_681 : entity work.gfmul
port map(
a=>a_3,
b=>"0100111001",
X=>mulr_3_681);

mulc_4_681 : entity work.gfmul
port map(
a=>a_4,
b=>"0010000001",
X=>mulr_4_681);

mulr_1_682<=a_1;
mulc_2_682 : entity work.gfmul
port map(
a=>a_2,
b=>"0011101100",
X=>mulr_2_682);

mulc_3_682 : entity work.gfmul
port map(
a=>a_3,
b=>"0011101101",
X=>mulr_3_682);

mulc_4_682 : entity work.gfmul
port map(
a=>a_4,
b=>"0000000001",
X=>mulr_4_682);

mulr_1_683<=a_1;
mulc_2_683 : entity work.gfmul
port map(
a=>a_2,
b=>"0111011000",
X=>mulr_2_683);

mulc_3_683 : entity work.gfmul
port map(
a=>a_3,
b=>"1110110100",
X=>mulr_3_683);

mulc_4_683 : entity work.gfmul
port map(
a=>a_4,
b=>"0000001000",
X=>mulr_4_683);

mulr_1_684<=a_1;
mulc_2_684 : entity work.gfmul
port map(
a=>a_2,
b=>"1110110000",
X=>mulr_2_684);

mulc_3_684 : entity work.gfmul
port map(
a=>a_3,
b=>"1011001011",
X=>mulr_3_684);

mulc_4_684 : entity work.gfmul
port map(
a=>a_4,
b=>"0001000000",
X=>mulr_4_684);

mulr_1_685<=a_1;
mulc_2_685 : entity work.gfmul
port map(
a=>a_2,
b=>"1101101001",
X=>mulr_2_685);

mulc_3_685 : entity work.gfmul
port map(
a=>a_3,
b=>"1100111110",
X=>mulr_3_685);

mulc_4_685 : entity work.gfmul
port map(
a=>a_4,
b=>"1000000000",
X=>mulr_4_685);

mulr_1_686<=a_1;
mulc_2_686 : entity work.gfmul
port map(
a=>a_2,
b=>"1011011011",
X=>mulr_2_686);

mulc_3_686 : entity work.gfmul
port map(
a=>a_3,
b=>"0011100011",
X=>mulr_3_686);

mulc_4_686 : entity work.gfmul
port map(
a=>a_4,
b=>"0000100100",
X=>mulr_4_686);

mulr_1_687<=a_1;
mulc_2_687 : entity work.gfmul
port map(
a=>a_2,
b=>"0110111111",
X=>mulr_2_687);

mulc_3_687 : entity work.gfmul
port map(
a=>a_3,
b=>"1110001100",
X=>mulr_3_687);

mulc_4_687 : entity work.gfmul
port map(
a=>a_4,
b=>"0100100000",
X=>mulr_4_687);

mulr_1_688<=a_1;
mulc_2_688 : entity work.gfmul
port map(
a=>a_2,
b=>"1101111110",
X=>mulr_2_688);

mulc_3_688 : entity work.gfmul
port map(
a=>a_3,
b=>"1000101011",
X=>mulr_3_688);

mulc_4_688 : entity work.gfmul
port map(
a=>a_4,
b=>"0100010010",
X=>mulr_4_688);

mulr_1_689<=a_1;
mulc_2_689 : entity work.gfmul
port map(
a=>a_2,
b=>"1011110101",
X=>mulr_2_689);

mulc_3_689 : entity work.gfmul
port map(
a=>a_3,
b=>"0010111110",
X=>mulr_3_689);

mulc_4_689 : entity work.gfmul
port map(
a=>a_4,
b=>"0010000010",
X=>mulr_4_689);

mulr_1_690<=a_1;
mulc_2_690 : entity work.gfmul
port map(
a=>a_2,
b=>"0111100011",
X=>mulr_2_690);

mulc_3_690 : entity work.gfmul
port map(
a=>a_3,
b=>"1011111000",
X=>mulr_3_690);

mulc_4_690 : entity work.gfmul
port map(
a=>a_4,
b=>"0000011001",
X=>mulr_4_690);

mulr_1_691<=a_1;
mulc_2_691 : entity work.gfmul
port map(
a=>a_2,
b=>"1111000110",
X=>mulr_2_691);

mulc_3_691 : entity work.gfmul
port map(
a=>a_3,
b=>"1111110010",
X=>mulr_3_691);

mulc_4_691 : entity work.gfmul
port map(
a=>a_4,
b=>"0011001000",
X=>mulr_4_691);

mulr_1_692<=a_1;
mulc_2_692 : entity work.gfmul
port map(
a=>a_2,
b=>"1110000101",
X=>mulr_2_692);

mulc_3_692 : entity work.gfmul
port map(
a=>a_3,
b=>"1111010011",
X=>mulr_3_692);

mulc_4_692 : entity work.gfmul
port map(
a=>a_4,
b=>"1001001001",
X=>mulr_4_692);

mulr_1_693<=a_1;
mulc_2_693 : entity work.gfmul
port map(
a=>a_2,
b=>"1100000011",
X=>mulr_2_693);

mulc_3_693 : entity work.gfmul
port map(
a=>a_3,
b=>"1101010111",
X=>mulr_3_693);

mulc_4_693 : entity work.gfmul
port map(
a=>a_4,
b=>"1001101100",
X=>mulr_4_693);

mulr_1_694<=a_1;
mulc_2_694 : entity work.gfmul
port map(
a=>a_2,
b=>"1000001111",
X=>mulr_2_694);

mulc_3_694 : entity work.gfmul
port map(
a=>a_3,
b=>"0101000111",
X=>mulr_3_694);

mulc_4_694 : entity work.gfmul
port map(
a=>a_4,
b=>"1101000100",
X=>mulr_4_694);

mulr_1_695<=a_1;
mulc_2_695 : entity work.gfmul
port map(
a=>a_2,
b=>"0000010111",
X=>mulr_2_695);

mulc_3_695 : entity work.gfmul
port map(
a=>a_3,
b=>"0100010101",
X=>mulr_3_695);

mulc_4_695 : entity work.gfmul
port map(
a=>a_4,
b=>"1000010110",
X=>mulr_4_695);

mulr_1_696<=a_1;
mulc_2_696 : entity work.gfmul
port map(
a=>a_2,
b=>"0000101110",
X=>mulr_2_696);

mulc_3_696 : entity work.gfmul
port map(
a=>a_3,
b=>"0001011101",
X=>mulr_3_696);

mulc_4_696 : entity work.gfmul
port map(
a=>a_4,
b=>"0010010100",
X=>mulr_4_696);

mulr_1_697<=a_1;
mulc_2_697 : entity work.gfmul
port map(
a=>a_2,
b=>"0001011100",
X=>mulr_2_697);

mulc_3_697 : entity work.gfmul
port map(
a=>a_3,
b=>"0101110100",
X=>mulr_3_697);

mulc_4_697 : entity work.gfmul
port map(
a=>a_4,
b=>"0010101001",
X=>mulr_4_697);

mulr_1_698<=a_1;
mulc_2_698 : entity work.gfmul
port map(
a=>a_2,
b=>"0010111000",
X=>mulr_2_698);

mulc_3_698 : entity work.gfmul
port map(
a=>a_3,
b=>"0111011001",
X=>mulr_3_698);

mulc_4_698 : entity work.gfmul
port map(
a=>a_4,
b=>"0101000001",
X=>mulr_4_698);

mulr_1_699<=a_1;
mulc_2_699 : entity work.gfmul
port map(
a=>a_2,
b=>"0101110000",
X=>mulr_2_699);

mulc_3_699 : entity work.gfmul
port map(
a=>a_3,
b=>"1101101101",
X=>mulr_3_699);

mulc_4_699 : entity work.gfmul
port map(
a=>a_4,
b=>"1000011010",
X=>mulr_4_699);

mulr_1_700<=a_1;
mulc_2_700 : entity work.gfmul
port map(
a=>a_2,
b=>"1011100000",
X=>mulr_2_700);

mulc_3_700 : entity work.gfmul
port map(
a=>a_3,
b=>"0110101111",
X=>mulr_3_700);

mulc_4_700 : entity work.gfmul
port map(
a=>a_4,
b=>"0011110100",
X=>mulr_4_700);

mulr_1_701<=a_1;
mulc_2_701 : entity work.gfmul
port map(
a=>a_2,
b=>"0111001001",
X=>mulr_2_701);

mulc_3_701 : entity work.gfmul
port map(
a=>a_3,
b=>"1010110101",
X=>mulr_3_701);

mulc_4_701 : entity work.gfmul
port map(
a=>a_4,
b=>"1110101001",
X=>mulr_4_701);

mulr_1_702<=a_1;
mulc_2_702 : entity work.gfmul
port map(
a=>a_2,
b=>"1110010010",
X=>mulr_2_702);

mulc_3_702 : entity work.gfmul
port map(
a=>a_3,
b=>"1011000110",
X=>mulr_3_702);

mulc_4_702 : entity work.gfmul
port map(
a=>a_4,
b=>"0101110111",
X=>mulr_4_702);

mulr_1_703<=a_1;
mulc_2_703 : entity work.gfmul
port map(
a=>a_2,
b=>"1100101101",
X=>mulr_2_703);

mulc_3_703 : entity work.gfmul
port map(
a=>a_3,
b=>"1100001010",
X=>mulr_3_703);

mulc_4_703 : entity work.gfmul
port map(
a=>a_4,
b=>"1110101010",
X=>mulr_4_703);

mulr_1_704<=a_1;
mulc_2_704 : entity work.gfmul
port map(
a=>a_2,
b=>"1001010011",
X=>mulr_2_704);

mulc_3_704 : entity work.gfmul
port map(
a=>a_3,
b=>"0000110011",
X=>mulr_3_704);

mulc_4_704 : entity work.gfmul
port map(
a=>a_4,
b=>"0101101111",
X=>mulr_4_704);

mulr_1_705<=a_1;
mulc_2_705 : entity work.gfmul
port map(
a=>a_2,
b=>"0010101111",
X=>mulr_2_705);

mulc_3_705 : entity work.gfmul
port map(
a=>a_3,
b=>"0011001100",
X=>mulr_3_705);

mulc_4_705 : entity work.gfmul
port map(
a=>a_4,
b=>"1101101010",
X=>mulr_4_705);

mulr_1_706<=a_1;
mulc_2_706 : entity work.gfmul
port map(
a=>a_2,
b=>"0101011110",
X=>mulr_2_706);

mulc_3_706 : entity work.gfmul
port map(
a=>a_3,
b=>"1100110000",
X=>mulr_3_706);

mulc_4_706 : entity work.gfmul
port map(
a=>a_4,
b=>"1101100110",
X=>mulr_4_706);

mulr_1_707<=a_1;
mulc_2_707 : entity work.gfmul
port map(
a=>a_2,
b=>"1010111100",
X=>mulr_2_707);

mulc_3_707 : entity work.gfmul
port map(
a=>a_3,
b=>"0011011011",
X=>mulr_3_707);

mulc_4_707 : entity work.gfmul
port map(
a=>a_4,
b=>"1100000110",
X=>mulr_4_707);

mulr_1_708<=a_1;
mulc_2_708 : entity work.gfmul
port map(
a=>a_2,
b=>"0101110001",
X=>mulr_2_708);

mulc_3_708 : entity work.gfmul
port map(
a=>a_3,
b=>"1101101100",
X=>mulr_3_708);

mulc_4_708 : entity work.gfmul
port map(
a=>a_4,
b=>"0000000110",
X=>mulr_4_708);

mulr_1_709<=a_1;
mulc_2_709 : entity work.gfmul
port map(
a=>a_2,
b=>"1011100010",
X=>mulr_2_709);

mulc_3_709 : entity work.gfmul
port map(
a=>a_3,
b=>"0110101011",
X=>mulr_3_709);

mulc_4_709 : entity work.gfmul
port map(
a=>a_4,
b=>"0000110000",
X=>mulr_4_709);

mulr_1_710<=a_1;
mulc_2_710 : entity work.gfmul
port map(
a=>a_2,
b=>"0111001101",
X=>mulr_2_710);

mulc_3_710 : entity work.gfmul
port map(
a=>a_3,
b=>"1010100101",
X=>mulr_3_710);

mulc_4_710 : entity work.gfmul
port map(
a=>a_4,
b=>"0110000000",
X=>mulr_4_710);

mulr_1_711<=a_1;
mulc_2_711 : entity work.gfmul
port map(
a=>a_2,
b=>"1110011010",
X=>mulr_2_711);

mulc_3_711 : entity work.gfmul
port map(
a=>a_3,
b=>"1010000110",
X=>mulr_3_711);

mulc_4_711 : entity work.gfmul
port map(
a=>a_4,
b=>"0000011011",
X=>mulr_4_711);

mulr_1_712<=a_1;
mulc_2_712 : entity work.gfmul
port map(
a=>a_2,
b=>"1100111101",
X=>mulr_2_712);

mulc_3_712 : entity work.gfmul
port map(
a=>a_3,
b=>"1000001010",
X=>mulr_3_712);

mulc_4_712 : entity work.gfmul
port map(
a=>a_4,
b=>"0011011000",
X=>mulr_4_712);

mulr_1_713<=a_1;
mulc_2_713 : entity work.gfmul
port map(
a=>a_2,
b=>"1001110011",
X=>mulr_2_713);

mulc_3_713 : entity work.gfmul
port map(
a=>a_3,
b=>"0000111010",
X=>mulr_3_713);

mulc_4_713 : entity work.gfmul
port map(
a=>a_4,
b=>"1011001001",
X=>mulr_4_713);

mulr_1_714<=a_1;
mulc_2_714 : entity work.gfmul
port map(
a=>a_2,
b=>"0011101111",
X=>mulr_2_714);

mulc_3_714 : entity work.gfmul
port map(
a=>a_3,
b=>"0011101000",
X=>mulr_3_714);

mulc_4_714 : entity work.gfmul
port map(
a=>a_4,
b=>"1001100101",
X=>mulr_4_714);

mulr_1_715<=a_1;
mulc_2_715 : entity work.gfmul
port map(
a=>a_2,
b=>"0111011110",
X=>mulr_2_715);

mulc_3_715 : entity work.gfmul
port map(
a=>a_3,
b=>"1110100000",
X=>mulr_3_715);

mulc_4_715 : entity work.gfmul
port map(
a=>a_4,
b=>"1100001100",
X=>mulr_4_715);

mulr_1_716<=a_1;
mulc_2_716 : entity work.gfmul
port map(
a=>a_2,
b=>"1110111100",
X=>mulr_2_716);

mulc_3_716 : entity work.gfmul
port map(
a=>a_3,
b=>"1010011011",
X=>mulr_3_716);

mulc_4_716 : entity work.gfmul
port map(
a=>a_4,
b=>"0001010110",
X=>mulr_4_716);

mulr_1_717<=a_1;
mulc_2_717 : entity work.gfmul
port map(
a=>a_2,
b=>"1101110001",
X=>mulr_2_717);

mulc_3_717 : entity work.gfmul
port map(
a=>a_3,
b=>"1001111110",
X=>mulr_3_717);

mulc_4_717 : entity work.gfmul
port map(
a=>a_4,
b=>"1010110000",
X=>mulr_4_717);

mulr_1_718<=a_1;
mulc_2_718 : entity work.gfmul
port map(
a=>a_2,
b=>"1011101011",
X=>mulr_2_718);

mulc_3_718 : entity work.gfmul
port map(
a=>a_3,
b=>"0111101010",
X=>mulr_3_718);

mulc_4_718 : entity work.gfmul
port map(
a=>a_4,
b=>"0110101101",
X=>mulr_4_718);

mulr_1_719<=a_1;
mulc_2_719 : entity work.gfmul
port map(
a=>a_2,
b=>"0111011111",
X=>mulr_2_719);

mulc_3_719 : entity work.gfmul
port map(
a=>a_3,
b=>"1110100001",
X=>mulr_3_719);

mulc_4_719 : entity work.gfmul
port map(
a=>a_4,
b=>"0101110011",
X=>mulr_4_719);

mulr_1_720<=a_1;
mulc_2_720 : entity work.gfmul
port map(
a=>a_2,
b=>"1110111110",
X=>mulr_2_720);

mulc_3_720 : entity work.gfmul
port map(
a=>a_3,
b=>"1010011111",
X=>mulr_3_720);

mulc_4_720 : entity work.gfmul
port map(
a=>a_4,
b=>"1110001010",
X=>mulr_4_720);

mulr_1_721<=a_1;
mulc_2_721 : entity work.gfmul
port map(
a=>a_2,
b=>"1101110101",
X=>mulr_2_721);

mulc_3_721 : entity work.gfmul
port map(
a=>a_3,
b=>"1001101110",
X=>mulr_3_721);

mulc_4_721 : entity work.gfmul
port map(
a=>a_4,
b=>"0001101111",
X=>mulr_4_721);

mulr_1_722<=a_1;
mulc_2_722 : entity work.gfmul
port map(
a=>a_2,
b=>"1011100011",
X=>mulr_2_722);

mulc_3_722 : entity work.gfmul
port map(
a=>a_3,
b=>"0110101010",
X=>mulr_3_722);

mulc_4_722 : entity work.gfmul
port map(
a=>a_4,
b=>"1101111000",
X=>mulr_4_722);

mulr_1_723<=a_1;
mulc_2_723 : entity work.gfmul
port map(
a=>a_2,
b=>"0111001111",
X=>mulr_2_723);

mulc_3_723 : entity work.gfmul
port map(
a=>a_3,
b=>"1010100001",
X=>mulr_3_723);

mulc_4_723 : entity work.gfmul
port map(
a=>a_4,
b=>"1111110110",
X=>mulr_4_723);

mulr_1_724<=a_1;
mulc_2_724 : entity work.gfmul
port map(
a=>a_2,
b=>"1110011110",
X=>mulr_2_724);

mulc_3_724 : entity work.gfmul
port map(
a=>a_3,
b=>"1010010110",
X=>mulr_3_724);

mulc_4_724 : entity work.gfmul
port map(
a=>a_4,
b=>"1110001111",
X=>mulr_4_724);

mulr_1_725<=a_1;
mulc_2_725 : entity work.gfmul
port map(
a=>a_2,
b=>"1100110101",
X=>mulr_2_725);

mulc_3_725 : entity work.gfmul
port map(
a=>a_3,
b=>"1001001010",
X=>mulr_3_725);

mulc_4_725 : entity work.gfmul
port map(
a=>a_4,
b=>"0001000111",
X=>mulr_4_725);

mulr_1_726<=a_1;
mulc_2_726 : entity work.gfmul
port map(
a=>a_2,
b=>"1001100011",
X=>mulr_2_726);

mulc_3_726 : entity work.gfmul
port map(
a=>a_3,
b=>"0100111010",
X=>mulr_3_726);

mulc_4_726 : entity work.gfmul
port map(
a=>a_4,
b=>"1000111000",
X=>mulr_4_726);

mulr_1_727<=a_1;
mulc_2_727 : entity work.gfmul
port map(
a=>a_2,
b=>"0011001111",
X=>mulr_2_727);

mulc_3_727 : entity work.gfmul
port map(
a=>a_3,
b=>"0011100001",
X=>mulr_3_727);

mulc_4_727 : entity work.gfmul
port map(
a=>a_4,
b=>"0111100100",
X=>mulr_4_727);

mulr_1_728<=a_1;
mulc_2_728 : entity work.gfmul
port map(
a=>a_2,
b=>"0110011110",
X=>mulr_2_728);

mulc_3_728 : entity work.gfmul
port map(
a=>a_3,
b=>"1110000100",
X=>mulr_3_728);

mulc_4_728 : entity work.gfmul
port map(
a=>a_4,
b=>"1100111011",
X=>mulr_4_728);

mulr_1_729<=a_1;
mulc_2_729 : entity work.gfmul
port map(
a=>a_2,
b=>"1100111100",
X=>mulr_2_729);

mulc_3_729 : entity work.gfmul
port map(
a=>a_3,
b=>"1000001011",
X=>mulr_3_729);

mulc_4_729 : entity work.gfmul
port map(
a=>a_4,
b=>"0111101110",
X=>mulr_4_729);

mulr_1_730<=a_1;
mulc_2_730 : entity work.gfmul
port map(
a=>a_2,
b=>"1001110001",
X=>mulr_2_730);

mulc_3_730 : entity work.gfmul
port map(
a=>a_3,
b=>"0000111110",
X=>mulr_3_730);

mulc_4_730 : entity work.gfmul
port map(
a=>a_4,
b=>"1101101011",
X=>mulr_4_730);

mulr_1_731<=a_1;
mulc_2_731 : entity work.gfmul
port map(
a=>a_2,
b=>"0011101011",
X=>mulr_2_731);

mulc_3_731 : entity work.gfmul
port map(
a=>a_3,
b=>"0011111000",
X=>mulr_3_731);

mulc_4_731 : entity work.gfmul
port map(
a=>a_4,
b=>"1101101110",
X=>mulr_4_731);

mulr_1_732<=a_1;
mulc_2_732 : entity work.gfmul
port map(
a=>a_2,
b=>"0111010110",
X=>mulr_2_732);

mulc_3_732 : entity work.gfmul
port map(
a=>a_3,
b=>"1111100000",
X=>mulr_3_732);

mulc_4_732 : entity work.gfmul
port map(
a=>a_4,
b=>"1101000110",
X=>mulr_4_732);

mulr_1_733<=a_1;
mulc_2_733 : entity work.gfmul
port map(
a=>a_2,
b=>"1110101100",
X=>mulr_2_733);

mulc_3_733 : entity work.gfmul
port map(
a=>a_3,
b=>"1110011011",
X=>mulr_3_733);

mulc_4_733 : entity work.gfmul
port map(
a=>a_4,
b=>"1000000110",
X=>mulr_4_733);

mulr_1_734<=a_1;
mulc_2_734 : entity work.gfmul
port map(
a=>a_2,
b=>"1101010001",
X=>mulr_2_734);

mulc_3_734 : entity work.gfmul
port map(
a=>a_3,
b=>"1001110111",
X=>mulr_3_734);

mulc_4_734 : entity work.gfmul
port map(
a=>a_4,
b=>"0000010100",
X=>mulr_4_734);

mulr_1_735<=a_1;
mulc_2_735 : entity work.gfmul
port map(
a=>a_2,
b=>"1010101011",
X=>mulr_2_735);

mulc_3_735 : entity work.gfmul
port map(
a=>a_3,
b=>"0111001110",
X=>mulr_3_735);

mulc_4_735 : entity work.gfmul
port map(
a=>a_4,
b=>"0010100000",
X=>mulr_4_735);

mulr_1_736<=a_1;
mulc_2_736 : entity work.gfmul
port map(
a=>a_2,
b=>"0101011111",
X=>mulr_2_736);

mulc_3_736 : entity work.gfmul
port map(
a=>a_3,
b=>"1100110001",
X=>mulr_3_736);

mulc_4_736 : entity work.gfmul
port map(
a=>a_4,
b=>"0100001001",
X=>mulr_4_736);

mulr_1_737<=a_1;
mulc_2_737 : entity work.gfmul
port map(
a=>a_2,
b=>"1010111110",
X=>mulr_2_737);

mulc_3_737 : entity work.gfmul
port map(
a=>a_3,
b=>"0011011111",
X=>mulr_3_737);

mulc_4_737 : entity work.gfmul
port map(
a=>a_4,
b=>"0001011010",
X=>mulr_4_737);

mulr_1_738<=a_1;
mulc_2_738 : entity work.gfmul
port map(
a=>a_2,
b=>"0101110101",
X=>mulr_2_738);

mulc_3_738 : entity work.gfmul
port map(
a=>a_3,
b=>"1101111100",
X=>mulr_3_738);

mulc_4_738 : entity work.gfmul
port map(
a=>a_4,
b=>"1011010000",
X=>mulr_4_738);

mulr_1_739<=a_1;
mulc_2_739 : entity work.gfmul
port map(
a=>a_2,
b=>"1011101010",
X=>mulr_2_739);

mulc_3_739 : entity work.gfmul
port map(
a=>a_3,
b=>"0111101011",
X=>mulr_3_739);

mulc_4_739 : entity work.gfmul
port map(
a=>a_4,
b=>"1010101101",
X=>mulr_4_739);

mulr_1_740<=a_1;
mulc_2_740 : entity work.gfmul
port map(
a=>a_2,
b=>"0111011101",
X=>mulr_2_740);

mulc_3_740 : entity work.gfmul
port map(
a=>a_3,
b=>"1110100101",
X=>mulr_3_740);

mulc_4_740 : entity work.gfmul
port map(
a=>a_4,
b=>"0101000101",
X=>mulr_4_740);

mulr_1_741<=a_1;
mulc_2_741 : entity work.gfmul
port map(
a=>a_2,
b=>"1110111010",
X=>mulr_2_741);

mulc_3_741 : entity work.gfmul
port map(
a=>a_3,
b=>"1010001111",
X=>mulr_3_741);

mulc_4_741 : entity work.gfmul
port map(
a=>a_4,
b=>"1000111010",
X=>mulr_4_741);

mulr_1_742<=a_1;
mulc_2_742 : entity work.gfmul
port map(
a=>a_2,
b=>"1101111101",
X=>mulr_2_742);

mulc_3_742 : entity work.gfmul
port map(
a=>a_3,
b=>"1000101110",
X=>mulr_3_742);

mulc_4_742 : entity work.gfmul
port map(
a=>a_4,
b=>"0111110100",
X=>mulr_4_742);

mulr_1_743<=a_1;
mulc_2_743 : entity work.gfmul
port map(
a=>a_2,
b=>"1011110011",
X=>mulr_2_743);

mulc_3_743 : entity work.gfmul
port map(
a=>a_3,
b=>"0010101010",
X=>mulr_3_743);

mulc_4_743 : entity work.gfmul
port map(
a=>a_4,
b=>"1110111011",
X=>mulr_4_743);

mulr_1_744<=a_1;
mulc_2_744 : entity work.gfmul
port map(
a=>a_2,
b=>"0111101111",
X=>mulr_2_744);

mulc_3_744 : entity work.gfmul
port map(
a=>a_3,
b=>"1010101000",
X=>mulr_3_744);

mulc_4_744 : entity work.gfmul
port map(
a=>a_4,
b=>"0111100111",
X=>mulr_4_744);

mulr_1_745<=a_1;
mulc_2_745 : entity work.gfmul
port map(
a=>a_2,
b=>"1111011110",
X=>mulr_2_745);

mulc_3_745 : entity work.gfmul
port map(
a=>a_3,
b=>"1010110010",
X=>mulr_3_745);

mulc_4_745 : entity work.gfmul
port map(
a=>a_4,
b=>"1100100011",
X=>mulr_4_745);

mulr_1_746<=a_1;
mulc_2_746 : entity work.gfmul
port map(
a=>a_2,
b=>"1110110101",
X=>mulr_2_746);

mulc_3_746 : entity work.gfmul
port map(
a=>a_3,
b=>"1011011010",
X=>mulr_3_746);

mulc_4_746 : entity work.gfmul
port map(
a=>a_4,
b=>"0100101110",
X=>mulr_4_746);

mulr_1_747<=a_1;
mulc_2_747 : entity work.gfmul
port map(
a=>a_2,
b=>"1101100011",
X=>mulr_2_747);

mulc_3_747 : entity work.gfmul
port map(
a=>a_3,
b=>"1101111010",
X=>mulr_3_747);

mulc_4_747 : entity work.gfmul
port map(
a=>a_4,
b=>"0101100010",
X=>mulr_4_747);

mulr_1_748<=a_1;
mulc_2_748 : entity work.gfmul
port map(
a=>a_2,
b=>"1011001111",
X=>mulr_2_748);

mulc_3_748 : entity work.gfmul
port map(
a=>a_3,
b=>"0111110011",
X=>mulr_3_748);

mulc_4_748 : entity work.gfmul
port map(
a=>a_4,
b=>"1100000010",
X=>mulr_4_748);

mulr_1_749<=a_1;
mulc_2_749 : entity work.gfmul
port map(
a=>a_2,
b=>"0110010111",
X=>mulr_2_749);

mulc_3_749 : entity work.gfmul
port map(
a=>a_3,
b=>"1111000101",
X=>mulr_3_749);

mulc_4_749 : entity work.gfmul
port map(
a=>a_4,
b=>"0000100110",
X=>mulr_4_749);

mulr_1_750<=a_1;
mulc_2_750 : entity work.gfmul
port map(
a=>a_2,
b=>"1100101110",
X=>mulr_2_750);

mulc_3_750 : entity work.gfmul
port map(
a=>a_3,
b=>"1100001111",
X=>mulr_3_750);

mulc_4_750 : entity work.gfmul
port map(
a=>a_4,
b=>"0100110000",
X=>mulr_4_750);

mulr_1_751<=a_1;
mulc_2_751 : entity work.gfmul
port map(
a=>a_2,
b=>"1001010101",
X=>mulr_2_751);

mulc_3_751 : entity work.gfmul
port map(
a=>a_3,
b=>"0000100111",
X=>mulr_3_751);

mulc_4_751 : entity work.gfmul
port map(
a=>a_4,
b=>"0110010010",
X=>mulr_4_751);

mulr_1_752<=a_1;
mulc_2_752 : entity work.gfmul
port map(
a=>a_2,
b=>"0010100011",
X=>mulr_2_752);

mulc_3_752 : entity work.gfmul
port map(
a=>a_3,
b=>"0010011100",
X=>mulr_3_752);

mulc_4_752 : entity work.gfmul
port map(
a=>a_4,
b=>"0010001011",
X=>mulr_4_752);

mulr_1_753<=a_1;
mulc_2_753 : entity work.gfmul
port map(
a=>a_2,
b=>"0101000110",
X=>mulr_2_753);

mulc_3_753 : entity work.gfmul
port map(
a=>a_3,
b=>"1001110000",
X=>mulr_3_753);

mulc_4_753 : entity work.gfmul
port map(
a=>a_4,
b=>"0001010001",
X=>mulr_4_753);

mulr_1_754<=a_1;
mulc_2_754 : entity work.gfmul
port map(
a=>a_2,
b=>"1010001100",
X=>mulr_2_754);

mulc_3_754 : entity work.gfmul
port map(
a=>a_3,
b=>"0111010010",
X=>mulr_3_754);

mulc_4_754 : entity work.gfmul
port map(
a=>a_4,
b=>"1010001000",
X=>mulr_4_754);

mulr_1_755<=a_1;
mulc_2_755 : entity work.gfmul
port map(
a=>a_2,
b=>"0100010001",
X=>mulr_2_755);

mulc_3_755 : entity work.gfmul
port map(
a=>a_3,
b=>"1101000001",
X=>mulr_3_755);

mulc_4_755 : entity work.gfmul
port map(
a=>a_4,
b=>"0001101101",
X=>mulr_4_755);

mulr_1_756<=a_1;
mulc_2_756 : entity work.gfmul
port map(
a=>a_2,
b=>"1000100010",
X=>mulr_2_756);

mulc_3_756 : entity work.gfmul
port map(
a=>a_3,
b=>"0100011111",
X=>mulr_3_756);

mulc_4_756 : entity work.gfmul
port map(
a=>a_4,
b=>"1101101000",
X=>mulr_4_756);

mulr_1_757<=a_1;
mulc_2_757 : entity work.gfmul
port map(
a=>a_2,
b=>"0001001101",
X=>mulr_2_757);

mulc_3_757 : entity work.gfmul
port map(
a=>a_3,
b=>"0001110101",
X=>mulr_3_757);

mulc_4_757 : entity work.gfmul
port map(
a=>a_4,
b=>"1101110110",
X=>mulr_4_757);

mulr_1_758<=a_1;
mulc_2_758 : entity work.gfmul
port map(
a=>a_2,
b=>"0010011010",
X=>mulr_2_758);

mulc_3_758 : entity work.gfmul
port map(
a=>a_3,
b=>"0111010100",
X=>mulr_3_758);

mulc_4_758 : entity work.gfmul
port map(
a=>a_4,
b=>"1110000110",
X=>mulr_4_758);

mulr_1_759<=a_1;
mulc_2_759 : entity work.gfmul
port map(
a=>a_2,
b=>"0100110100",
X=>mulr_2_759);

mulc_3_759 : entity work.gfmul
port map(
a=>a_3,
b=>"1101011001",
X=>mulr_3_759);

mulc_4_759 : entity work.gfmul
port map(
a=>a_4,
b=>"0000001111",
X=>mulr_4_759);

mulr_1_760<=a_1;
mulc_2_760 : entity work.gfmul
port map(
a=>a_2,
b=>"1001101000",
X=>mulr_2_760);

mulc_3_760 : entity work.gfmul
port map(
a=>a_3,
b=>"0101111111",
X=>mulr_3_760);

mulc_4_760 : entity work.gfmul
port map(
a=>a_4,
b=>"0001111000",
X=>mulr_4_760);

mulr_1_761<=a_1;
mulc_2_761 : entity work.gfmul
port map(
a=>a_2,
b=>"0011011001",
X=>mulr_2_761);

mulc_3_761 : entity work.gfmul
port map(
a=>a_3,
b=>"0111110101",
X=>mulr_3_761);

mulc_4_761 : entity work.gfmul
port map(
a=>a_4,
b=>"1111000000",
X=>mulr_4_761);

mulr_1_762<=a_1;
mulc_2_762 : entity work.gfmul
port map(
a=>a_2,
b=>"0110110010",
X=>mulr_2_762);

mulc_3_762 : entity work.gfmul
port map(
a=>a_3,
b=>"1111011101",
X=>mulr_3_762);

mulc_4_762 : entity work.gfmul
port map(
a=>a_4,
b=>"1000111111",
X=>mulr_4_762);

mulr_1_763<=a_1;
mulc_2_763 : entity work.gfmul
port map(
a=>a_2,
b=>"1101100100",
X=>mulr_2_763);

mulc_3_763 : entity work.gfmul
port map(
a=>a_3,
b=>"1101101111",
X=>mulr_3_763);

mulc_4_763 : entity work.gfmul
port map(
a=>a_4,
b=>"0111011100",
X=>mulr_4_763);

mulr_1_764<=a_1;
mulc_2_764 : entity work.gfmul
port map(
a=>a_2,
b=>"1011000001",
X=>mulr_2_764);

mulc_3_764 : entity work.gfmul
port map(
a=>a_3,
b=>"0110100111",
X=>mulr_3_764);

mulc_4_764 : entity work.gfmul
port map(
a=>a_4,
b=>"1011111011",
X=>mulr_4_764);

mulr_1_765<=a_1;
mulc_2_765 : entity work.gfmul
port map(
a=>a_2,
b=>"0110001011",
X=>mulr_2_765);

mulc_3_765 : entity work.gfmul
port map(
a=>a_3,
b=>"1010010101",
X=>mulr_3_765);

mulc_4_765 : entity work.gfmul
port map(
a=>a_4,
b=>"1111110101",
X=>mulr_4_765);

mulr_1_766<=a_1;
mulc_2_766 : entity work.gfmul
port map(
a=>a_2,
b=>"1100010110",
X=>mulr_2_766);

mulc_3_766 : entity work.gfmul
port map(
a=>a_3,
b=>"1001000110",
X=>mulr_3_766);

mulc_4_766 : entity work.gfmul
port map(
a=>a_4,
b=>"1110010111",
X=>mulr_4_766);

mulr_1_767<=a_1;
mulc_2_767 : entity work.gfmul
port map(
a=>a_2,
b=>"1000100101",
X=>mulr_2_767);

mulc_3_767 : entity work.gfmul
port map(
a=>a_3,
b=>"0100001010",
X=>mulr_3_767);

mulc_4_767 : entity work.gfmul
port map(
a=>a_4,
b=>"0010000111",
X=>mulr_4_767);

mulr_1_768<=a_1;
mulc_2_768 : entity work.gfmul
port map(
a=>a_2,
b=>"0001000011",
X=>mulr_2_768);

mulc_3_768 : entity work.gfmul
port map(
a=>a_3,
b=>"0000100001",
X=>mulr_3_768);

mulc_4_768 : entity work.gfmul
port map(
a=>a_4,
b=>"0000110001",
X=>mulr_4_768);

mulr_1_769<=a_1;
mulc_2_769 : entity work.gfmul
port map(
a=>a_2,
b=>"0010000110",
X=>mulr_2_769);

mulc_3_769 : entity work.gfmul
port map(
a=>a_3,
b=>"0010000100",
X=>mulr_3_769);

mulc_4_769 : entity work.gfmul
port map(
a=>a_4,
b=>"0110001000",
X=>mulr_4_769);

mulr_1_770<=a_1;
mulc_2_770 : entity work.gfmul
port map(
a=>a_2,
b=>"0100001100",
X=>mulr_2_770);

mulc_3_770 : entity work.gfmul
port map(
a=>a_3,
b=>"1000010000",
X=>mulr_3_770);

mulc_4_770 : entity work.gfmul
port map(
a=>a_4,
b=>"0001011011",
X=>mulr_4_770);

mulr_1_771<=a_1;
mulc_2_771 : entity work.gfmul
port map(
a=>a_2,
b=>"1000011000",
X=>mulr_2_771);

mulc_3_771 : entity work.gfmul
port map(
a=>a_3,
b=>"0001010010",
X=>mulr_3_771);

mulc_4_771 : entity work.gfmul
port map(
a=>a_4,
b=>"1011011000",
X=>mulr_4_771);

mulr_1_772<=a_1;
mulc_2_772 : entity work.gfmul
port map(
a=>a_2,
b=>"0000111001",
X=>mulr_2_772);

mulc_3_772 : entity work.gfmul
port map(
a=>a_3,
b=>"0101001000",
X=>mulr_3_772);

mulc_4_772 : entity work.gfmul
port map(
a=>a_4,
b=>"1011101101",
X=>mulr_4_772);

mulr_1_773<=a_1;
mulc_2_773 : entity work.gfmul
port map(
a=>a_2,
b=>"0001110010",
X=>mulr_2_773);

mulc_3_773 : entity work.gfmul
port map(
a=>a_3,
b=>"0100101001",
X=>mulr_3_773);

mulc_4_773 : entity work.gfmul
port map(
a=>a_4,
b=>"1101000101",
X=>mulr_4_773);

mulr_1_774<=a_1;
mulc_2_774 : entity work.gfmul
port map(
a=>a_2,
b=>"0011100100",
X=>mulr_2_774);

mulc_3_774 : entity work.gfmul
port map(
a=>a_3,
b=>"0010101101",
X=>mulr_3_774);

mulc_4_774 : entity work.gfmul
port map(
a=>a_4,
b=>"1000011110",
X=>mulr_4_774);

mulr_1_775<=a_1;
mulc_2_775 : entity work.gfmul
port map(
a=>a_2,
b=>"0111001000",
X=>mulr_2_775);

mulc_3_775 : entity work.gfmul
port map(
a=>a_3,
b=>"1010110100",
X=>mulr_3_775);

mulc_4_775 : entity work.gfmul
port map(
a=>a_4,
b=>"0011010100",
X=>mulr_4_775);

mulr_1_776<=a_1;
mulc_2_776 : entity work.gfmul
port map(
a=>a_2,
b=>"1110010000",
X=>mulr_2_776);

mulc_3_776 : entity work.gfmul
port map(
a=>a_3,
b=>"1011000010",
X=>mulr_3_776);

mulc_4_776 : entity work.gfmul
port map(
a=>a_4,
b=>"1010101001",
X=>mulr_4_776);

mulr_1_777<=a_1;
mulc_2_777 : entity work.gfmul
port map(
a=>a_2,
b=>"1100101001",
X=>mulr_2_777);

mulc_3_777 : entity work.gfmul
port map(
a=>a_3,
b=>"1100011010",
X=>mulr_3_777);

mulc_4_777 : entity work.gfmul
port map(
a=>a_4,
b=>"0101100101",
X=>mulr_4_777);

mulr_1_778<=a_1;
mulc_2_778 : entity work.gfmul
port map(
a=>a_2,
b=>"1001011011",
X=>mulr_2_778);

mulc_3_778 : entity work.gfmul
port map(
a=>a_3,
b=>"0001110011",
X=>mulr_3_778);

mulc_4_778 : entity work.gfmul
port map(
a=>a_4,
b=>"1100111010",
X=>mulr_4_778);

mulr_1_779<=a_1;
mulc_2_779 : entity work.gfmul
port map(
a=>a_2,
b=>"0010111111",
X=>mulr_2_779);

mulc_3_779 : entity work.gfmul
port map(
a=>a_3,
b=>"0111001100",
X=>mulr_3_779);

mulc_4_779 : entity work.gfmul
port map(
a=>a_4,
b=>"0111100110",
X=>mulr_4_779);

mulr_1_780<=a_1;
mulc_2_780 : entity work.gfmul
port map(
a=>a_2,
b=>"0101111110",
X=>mulr_2_780);

mulc_3_780 : entity work.gfmul
port map(
a=>a_3,
b=>"1100111001",
X=>mulr_3_780);

mulc_4_780 : entity work.gfmul
port map(
a=>a_4,
b=>"1100101011",
X=>mulr_4_780);

mulr_1_781<=a_1;
mulc_2_781 : entity work.gfmul
port map(
a=>a_2,
b=>"1011111100",
X=>mulr_2_781);

mulc_3_781 : entity work.gfmul
port map(
a=>a_3,
b=>"0011111111",
X=>mulr_3_781);

mulc_4_781 : entity work.gfmul
port map(
a=>a_4,
b=>"0101101110",
X=>mulr_4_781);

mulr_1_782<=a_1;
mulc_2_782 : entity work.gfmul
port map(
a=>a_2,
b=>"0111110001",
X=>mulr_2_782);

mulc_3_782 : entity work.gfmul
port map(
a=>a_3,
b=>"1111111100",
X=>mulr_3_782);

mulc_4_782 : entity work.gfmul
port map(
a=>a_4,
b=>"1101100010",
X=>mulr_4_782);

mulr_1_783<=a_1;
mulc_2_783 : entity work.gfmul
port map(
a=>a_2,
b=>"1111100010",
X=>mulr_2_783);

mulc_3_783 : entity work.gfmul
port map(
a=>a_3,
b=>"1111101011",
X=>mulr_3_783);

mulc_4_783 : entity work.gfmul
port map(
a=>a_4,
b=>"1100100110",
X=>mulr_4_783);

mulr_1_784<=a_1;
mulc_2_784 : entity work.gfmul
port map(
a=>a_2,
b=>"1111001101",
X=>mulr_2_784);

mulc_3_784 : entity work.gfmul
port map(
a=>a_3,
b=>"1110110111",
X=>mulr_3_784);

mulc_4_784 : entity work.gfmul
port map(
a=>a_4,
b=>"0100000110",
X=>mulr_4_784);

mulr_1_785<=a_1;
mulc_2_785 : entity work.gfmul
port map(
a=>a_2,
b=>"1110010011",
X=>mulr_2_785);

mulc_3_785 : entity work.gfmul
port map(
a=>a_3,
b=>"1011000111",
X=>mulr_3_785);

mulc_4_785 : entity work.gfmul
port map(
a=>a_4,
b=>"0000100010",
X=>mulr_4_785);

mulr_1_786<=a_1;
mulc_2_786 : entity work.gfmul
port map(
a=>a_2,
b=>"1100101111",
X=>mulr_2_786);

mulc_3_786 : entity work.gfmul
port map(
a=>a_3,
b=>"1100001110",
X=>mulr_3_786);

mulc_4_786 : entity work.gfmul
port map(
a=>a_4,
b=>"0100010000",
X=>mulr_4_786);

mulr_1_787<=a_1;
mulc_2_787 : entity work.gfmul
port map(
a=>a_2,
b=>"1001010111",
X=>mulr_2_787);

mulc_3_787 : entity work.gfmul
port map(
a=>a_3,
b=>"0000100011",
X=>mulr_3_787);

mulc_4_787 : entity work.gfmul
port map(
a=>a_4,
b=>"0010010010",
X=>mulr_4_787);

mulr_1_788<=a_1;
mulc_2_788 : entity work.gfmul
port map(
a=>a_2,
b=>"0010100111",
X=>mulr_2_788);

mulc_3_788 : entity work.gfmul
port map(
a=>a_3,
b=>"0010001100",
X=>mulr_3_788);

mulc_4_788 : entity work.gfmul
port map(
a=>a_4,
b=>"0010011001",
X=>mulr_4_788);

mulr_1_789<=a_1;
mulc_2_789 : entity work.gfmul
port map(
a=>a_2,
b=>"0101001110",
X=>mulr_2_789);

mulc_3_789 : entity work.gfmul
port map(
a=>a_3,
b=>"1000110000",
X=>mulr_3_789);

mulc_4_789 : entity work.gfmul
port map(
a=>a_4,
b=>"0011000001",
X=>mulr_4_789);

mulr_1_790<=a_1;
mulc_2_790 : entity work.gfmul
port map(
a=>a_2,
b=>"1010011100",
X=>mulr_2_790);

mulc_3_790 : entity work.gfmul
port map(
a=>a_3,
b=>"0011010010",
X=>mulr_3_790);

mulc_4_790 : entity work.gfmul
port map(
a=>a_4,
b=>"1000000001",
X=>mulr_4_790);

mulr_1_791<=a_1;
mulc_2_791 : entity work.gfmul
port map(
a=>a_2,
b=>"0100110001",
X=>mulr_2_791);

mulc_3_791 : entity work.gfmul
port map(
a=>a_3,
b=>"1101001000",
X=>mulr_3_791);

mulc_4_791 : entity work.gfmul
port map(
a=>a_4,
b=>"0000101100",
X=>mulr_4_791);

mulr_1_792<=a_1;
mulc_2_792 : entity work.gfmul
port map(
a=>a_2,
b=>"1001100010",
X=>mulr_2_792);

mulc_3_792 : entity work.gfmul
port map(
a=>a_3,
b=>"0100111011",
X=>mulr_3_792);

mulc_4_792 : entity work.gfmul
port map(
a=>a_4,
b=>"0101100000",
X=>mulr_4_792);

mulr_1_793<=a_1;
mulc_2_793 : entity work.gfmul
port map(
a=>a_2,
b=>"0011001101",
X=>mulr_2_793);

mulc_3_793 : entity work.gfmul
port map(
a=>a_3,
b=>"0011100101",
X=>mulr_3_793);

mulc_4_793 : entity work.gfmul
port map(
a=>a_4,
b=>"1100010010",
X=>mulr_4_793);

mulr_1_794<=a_1;
mulc_2_794 : entity work.gfmul
port map(
a=>a_2,
b=>"0110011010",
X=>mulr_2_794);

mulc_3_794 : entity work.gfmul
port map(
a=>a_3,
b=>"1110010100",
X=>mulr_3_794);

mulc_4_794 : entity work.gfmul
port map(
a=>a_4,
b=>"0010100110",
X=>mulr_4_794);

mulr_1_795<=a_1;
mulc_2_795 : entity work.gfmul
port map(
a=>a_2,
b=>"1100110100",
X=>mulr_2_795);

mulc_3_795 : entity work.gfmul
port map(
a=>a_3,
b=>"1001001011",
X=>mulr_3_795);

mulc_4_795 : entity work.gfmul
port map(
a=>a_4,
b=>"0100111001",
X=>mulr_4_795);

mulr_1_796<=a_1;
mulc_2_796 : entity work.gfmul
port map(
a=>a_2,
b=>"1001100001",
X=>mulr_2_796);

mulc_3_796 : entity work.gfmul
port map(
a=>a_3,
b=>"0100111110",
X=>mulr_3_796);

mulc_4_796 : entity work.gfmul
port map(
a=>a_4,
b=>"0111011010",
X=>mulr_4_796);

mulr_1_797<=a_1;
mulc_2_797 : entity work.gfmul
port map(
a=>a_2,
b=>"0011001011",
X=>mulr_2_797);

mulc_3_797 : entity work.gfmul
port map(
a=>a_3,
b=>"0011110001",
X=>mulr_3_797);

mulc_4_797 : entity work.gfmul
port map(
a=>a_4,
b=>"1011001011",
X=>mulr_4_797);

mulr_1_798<=a_1;
mulc_2_798 : entity work.gfmul
port map(
a=>a_2,
b=>"0110010110",
X=>mulr_2_798);

mulc_3_798 : entity work.gfmul
port map(
a=>a_3,
b=>"1111000100",
X=>mulr_3_798);

mulc_4_798 : entity work.gfmul
port map(
a=>a_4,
b=>"1001110101",
X=>mulr_4_798);

mulr_1_799<=a_1;
mulc_2_799 : entity work.gfmul
port map(
a=>a_2,
b=>"1100101100",
X=>mulr_2_799);

mulc_3_799 : entity work.gfmul
port map(
a=>a_3,
b=>"1100001011",
X=>mulr_3_799);

mulc_4_799 : entity work.gfmul
port map(
a=>a_4,
b=>"1110001100",
X=>mulr_4_799);

mulr_1_800<=a_1;
mulc_2_800 : entity work.gfmul
port map(
a=>a_2,
b=>"1001010001",
X=>mulr_2_800);

mulc_3_800 : entity work.gfmul
port map(
a=>a_3,
b=>"0000110111",
X=>mulr_3_800);

mulc_4_800 : entity work.gfmul
port map(
a=>a_4,
b=>"0001011111",
X=>mulr_4_800);

mulr_1_801<=a_1;
mulc_2_801 : entity work.gfmul
port map(
a=>a_2,
b=>"0010101011",
X=>mulr_2_801);

mulc_3_801 : entity work.gfmul
port map(
a=>a_3,
b=>"0011011100",
X=>mulr_3_801);

mulc_4_801 : entity work.gfmul
port map(
a=>a_4,
b=>"1011111000",
X=>mulr_4_801);

mulr_1_802<=a_1;
mulc_2_802 : entity work.gfmul
port map(
a=>a_2,
b=>"0101010110",
X=>mulr_2_802);

mulc_3_802 : entity work.gfmul
port map(
a=>a_3,
b=>"1101110000",
X=>mulr_3_802);

mulc_4_802 : entity work.gfmul
port map(
a=>a_4,
b=>"1111101101",
X=>mulr_4_802);

mulr_1_803<=a_1;
mulc_2_803 : entity work.gfmul
port map(
a=>a_2,
b=>"1010101100",
X=>mulr_2_803);

mulc_3_803 : entity work.gfmul
port map(
a=>a_3,
b=>"0111011011",
X=>mulr_3_803);

mulc_4_803 : entity work.gfmul
port map(
a=>a_4,
b=>"1101010111",
X=>mulr_4_803);

mulr_1_804<=a_1;
mulc_2_804 : entity work.gfmul
port map(
a=>a_2,
b=>"0101010001",
X=>mulr_2_804);

mulc_3_804 : entity work.gfmul
port map(
a=>a_3,
b=>"1101100101",
X=>mulr_3_804);

mulc_4_804 : entity work.gfmul
port map(
a=>a_4,
b=>"1010001110",
X=>mulr_4_804);

mulr_1_805<=a_1;
mulc_2_805 : entity work.gfmul
port map(
a=>a_2,
b=>"1010100010",
X=>mulr_2_805);

mulc_3_805 : entity work.gfmul
port map(
a=>a_3,
b=>"0110001111",
X=>mulr_3_805);

mulc_4_805 : entity work.gfmul
port map(
a=>a_4,
b=>"0001011101",
X=>mulr_4_805);

mulr_1_806<=a_1;
mulc_2_806 : entity work.gfmul
port map(
a=>a_2,
b=>"0101001101",
X=>mulr_2_806);

mulc_3_806 : entity work.gfmul
port map(
a=>a_3,
b=>"1000110101",
X=>mulr_3_806);

mulc_4_806 : entity work.gfmul
port map(
a=>a_4,
b=>"1011101000",
X=>mulr_4_806);

mulr_1_807<=a_1;
mulc_2_807 : entity work.gfmul
port map(
a=>a_2,
b=>"1010011010",
X=>mulr_2_807);

mulc_3_807 : entity work.gfmul
port map(
a=>a_3,
b=>"0011000110",
X=>mulr_3_807);

mulc_4_807 : entity work.gfmul
port map(
a=>a_4,
b=>"1101101101",
X=>mulr_4_807);

mulr_1_808<=a_1;
mulc_2_808 : entity work.gfmul
port map(
a=>a_2,
b=>"0100111101",
X=>mulr_2_808);

mulc_3_808 : entity work.gfmul
port map(
a=>a_3,
b=>"1100011000",
X=>mulr_3_808);

mulc_4_808 : entity work.gfmul
port map(
a=>a_4,
b=>"1101011110",
X=>mulr_4_808);

mulr_1_809<=a_1;
mulc_2_809 : entity work.gfmul
port map(
a=>a_2,
b=>"1001111010",
X=>mulr_2_809);

mulc_3_809 : entity work.gfmul
port map(
a=>a_3,
b=>"0001111011",
X=>mulr_3_809);

mulc_4_809 : entity work.gfmul
port map(
a=>a_4,
b=>"1011000110",
X=>mulr_4_809);

mulr_1_810<=a_1;
mulc_2_810 : entity work.gfmul
port map(
a=>a_2,
b=>"0011111101",
X=>mulr_2_810);

mulc_3_810 : entity work.gfmul
port map(
a=>a_3,
b=>"0111101100",
X=>mulr_3_810);

mulc_4_810 : entity work.gfmul
port map(
a=>a_4,
b=>"1000011101",
X=>mulr_4_810);

mulr_1_811<=a_1;
mulc_2_811 : entity work.gfmul
port map(
a=>a_2,
b=>"0111111010",
X=>mulr_2_811);

mulc_3_811 : entity work.gfmul
port map(
a=>a_3,
b=>"1110111001",
X=>mulr_3_811);

mulc_4_811 : entity work.gfmul
port map(
a=>a_4,
b=>"0011001100",
X=>mulr_4_811);

mulr_1_812<=a_1;
mulc_2_812 : entity work.gfmul
port map(
a=>a_2,
b=>"1111110100",
X=>mulr_2_812);

mulc_3_812 : entity work.gfmul
port map(
a=>a_3,
b=>"1011111111",
X=>mulr_3_812);

mulc_4_812 : entity work.gfmul
port map(
a=>a_4,
b=>"1001101001",
X=>mulr_4_812);

mulr_1_813<=a_1;
mulc_2_813 : entity work.gfmul
port map(
a=>a_2,
b=>"1111100001",
X=>mulr_2_813);

mulc_3_813 : entity work.gfmul
port map(
a=>a_3,
b=>"1111101110",
X=>mulr_3_813);

mulc_4_813 : entity work.gfmul
port map(
a=>a_4,
b=>"1101101100",
X=>mulr_4_813);

mulr_1_814<=a_1;
mulc_2_814 : entity work.gfmul
port map(
a=>a_2,
b=>"1111001011",
X=>mulr_2_814);

mulc_3_814 : entity work.gfmul
port map(
a=>a_3,
b=>"1110100011",
X=>mulr_3_814);

mulc_4_814 : entity work.gfmul
port map(
a=>a_4,
b=>"1101010110",
X=>mulr_4_814);

mulr_1_815<=a_1;
mulc_2_815 : entity work.gfmul
port map(
a=>a_2,
b=>"1110011111",
X=>mulr_2_815);

mulc_3_815 : entity work.gfmul
port map(
a=>a_3,
b=>"1010010111",
X=>mulr_3_815);

mulc_4_815 : entity work.gfmul
port map(
a=>a_4,
b=>"1010000110",
X=>mulr_4_815);

mulr_1_816<=a_1;
mulc_2_816 : entity work.gfmul
port map(
a=>a_2,
b=>"1100110111",
X=>mulr_2_816);

mulc_3_816 : entity work.gfmul
port map(
a=>a_3,
b=>"1001001110",
X=>mulr_3_816);

mulc_4_816 : entity work.gfmul
port map(
a=>a_4,
b=>"0000011101",
X=>mulr_4_816);

mulr_1_817<=a_1;
mulc_2_817 : entity work.gfmul
port map(
a=>a_2,
b=>"1001100111",
X=>mulr_2_817);

mulc_3_817 : entity work.gfmul
port map(
a=>a_3,
b=>"0100101010",
X=>mulr_3_817);

mulc_4_817 : entity work.gfmul
port map(
a=>a_4,
b=>"0011101000",
X=>mulr_4_817);

mulr_1_818<=a_1;
mulc_2_818 : entity work.gfmul
port map(
a=>a_2,
b=>"0011000111",
X=>mulr_2_818);

mulc_3_818 : entity work.gfmul
port map(
a=>a_3,
b=>"0010100001",
X=>mulr_3_818);

mulc_4_818 : entity work.gfmul
port map(
a=>a_4,
b=>"1101001001",
X=>mulr_4_818);

mulr_1_819<=a_1;
mulc_2_819 : entity work.gfmul
port map(
a=>a_2,
b=>"0110001110",
X=>mulr_2_819);

mulc_3_819 : entity work.gfmul
port map(
a=>a_3,
b=>"1010000100",
X=>mulr_3_819);

mulc_4_819 : entity work.gfmul
port map(
a=>a_4,
b=>"1001111110",
X=>mulr_4_819);

mulr_1_820<=a_1;
mulc_2_820 : entity work.gfmul
port map(
a=>a_2,
b=>"1100011100",
X=>mulr_2_820);

mulc_3_820 : entity work.gfmul
port map(
a=>a_3,
b=>"1000000010",
X=>mulr_3_820);

mulc_4_820 : entity work.gfmul
port map(
a=>a_4,
b=>"1111010100",
X=>mulr_4_820);

mulr_1_821<=a_1;
mulc_2_821 : entity work.gfmul
port map(
a=>a_2,
b=>"1000110001",
X=>mulr_2_821);

mulc_3_821 : entity work.gfmul
port map(
a=>a_3,
b=>"0000011010",
X=>mulr_3_821);

mulc_4_821 : entity work.gfmul
port map(
a=>a_4,
b=>"1010011111",
X=>mulr_4_821);

mulr_1_822<=a_1;
mulc_2_822 : entity work.gfmul
port map(
a=>a_2,
b=>"0001101011",
X=>mulr_2_822);

mulc_3_822 : entity work.gfmul
port map(
a=>a_3,
b=>"0001101000",
X=>mulr_3_822);

mulc_4_822 : entity work.gfmul
port map(
a=>a_4,
b=>"0011010101",
X=>mulr_4_822);

mulr_1_823<=a_1;
mulc_2_823 : entity work.gfmul
port map(
a=>a_2,
b=>"0011010110",
X=>mulr_2_823);

mulc_3_823 : entity work.gfmul
port map(
a=>a_3,
b=>"0110100000",
X=>mulr_3_823);

mulc_4_823 : entity work.gfmul
port map(
a=>a_4,
b=>"1010100001",
X=>mulr_4_823);

mulr_1_824<=a_1;
mulc_2_824 : entity work.gfmul
port map(
a=>a_2,
b=>"0110101100",
X=>mulr_2_824);

mulc_3_824 : entity work.gfmul
port map(
a=>a_3,
b=>"1010001001",
X=>mulr_3_824);

mulc_4_824 : entity work.gfmul
port map(
a=>a_4,
b=>"0100100101",
X=>mulr_4_824);

mulr_1_825<=a_1;
mulc_2_825 : entity work.gfmul
port map(
a=>a_2,
b=>"1101011000",
X=>mulr_2_825);

mulc_3_825 : entity work.gfmul
port map(
a=>a_3,
b=>"1000110110",
X=>mulr_3_825);

mulc_4_825 : entity work.gfmul
port map(
a=>a_4,
b=>"0100111010",
X=>mulr_4_825);

mulr_1_826<=a_1;
mulc_2_826 : entity work.gfmul
port map(
a=>a_2,
b=>"1010111001",
X=>mulr_2_826);

mulc_3_826 : entity work.gfmul
port map(
a=>a_3,
b=>"0011001010",
X=>mulr_3_826);

mulc_4_826 : entity work.gfmul
port map(
a=>a_4,
b=>"0111000010",
X=>mulr_4_826);

mulr_1_827<=a_1;
mulc_2_827 : entity work.gfmul
port map(
a=>a_2,
b=>"0101111011",
X=>mulr_2_827);

mulc_3_827 : entity work.gfmul
port map(
a=>a_3,
b=>"1100101000",
X=>mulr_3_827);

mulc_4_827 : entity work.gfmul
port map(
a=>a_4,
b=>"1000001011",
X=>mulr_4_827);

mulr_1_828<=a_1;
mulc_2_828 : entity work.gfmul
port map(
a=>a_2,
b=>"1011110110",
X=>mulr_2_828);

mulc_3_828 : entity work.gfmul
port map(
a=>a_3,
b=>"0010111011",
X=>mulr_3_828);

mulc_4_828 : entity work.gfmul
port map(
a=>a_4,
b=>"0001111100",
X=>mulr_4_828);

mulr_1_829<=a_1;
mulc_2_829 : entity work.gfmul
port map(
a=>a_2,
b=>"0111100101",
X=>mulr_2_829);

mulc_3_829 : entity work.gfmul
port map(
a=>a_3,
b=>"1011101100",
X=>mulr_3_829);

mulc_4_829 : entity work.gfmul
port map(
a=>a_4,
b=>"1111100000",
X=>mulr_4_829);

mulr_1_830<=a_1;
mulc_2_830 : entity work.gfmul
port map(
a=>a_2,
b=>"1111001010",
X=>mulr_2_830);

mulc_3_830 : entity work.gfmul
port map(
a=>a_3,
b=>"1110100010",
X=>mulr_3_830);

mulc_4_830 : entity work.gfmul
port map(
a=>a_4,
b=>"1100111111",
X=>mulr_4_830);

mulr_1_831<=a_1;
mulc_2_831 : entity work.gfmul
port map(
a=>a_2,
b=>"1110011101",
X=>mulr_2_831);

mulc_3_831 : entity work.gfmul
port map(
a=>a_3,
b=>"1010010011",
X=>mulr_3_831);

mulc_4_831 : entity work.gfmul
port map(
a=>a_4,
b=>"0111001110",
X=>mulr_4_831);

mulr_1_832<=a_1;
mulc_2_832 : entity work.gfmul
port map(
a=>a_2,
b=>"1100110011",
X=>mulr_2_832);

mulc_3_832 : entity work.gfmul
port map(
a=>a_3,
b=>"1001011110",
X=>mulr_3_832);

mulc_4_832 : entity work.gfmul
port map(
a=>a_4,
b=>"1001101011",
X=>mulr_4_832);

mulr_1_833<=a_1;
mulc_2_833 : entity work.gfmul
port map(
a=>a_2,
b=>"1001101111",
X=>mulr_2_833);

mulc_3_833 : entity work.gfmul
port map(
a=>a_3,
b=>"0101101010",
X=>mulr_3_833);

mulc_4_833 : entity work.gfmul
port map(
a=>a_4,
b=>"1101111100",
X=>mulr_4_833);

mulr_1_834<=a_1;
mulc_2_834 : entity work.gfmul
port map(
a=>a_2,
b=>"0011010111",
X=>mulr_2_834);

mulc_3_834 : entity work.gfmul
port map(
a=>a_3,
b=>"0110100001",
X=>mulr_3_834);

mulc_4_834 : entity work.gfmul
port map(
a=>a_4,
b=>"1111010110",
X=>mulr_4_834);

mulr_1_835<=a_1;
mulc_2_835 : entity work.gfmul
port map(
a=>a_2,
b=>"0110101110",
X=>mulr_2_835);

mulc_3_835 : entity work.gfmul
port map(
a=>a_3,
b=>"1010001101",
X=>mulr_3_835);

mulc_4_835 : entity work.gfmul
port map(
a=>a_4,
b=>"1010001111",
X=>mulr_4_835);

mulr_1_836<=a_1;
mulc_2_836 : entity work.gfmul
port map(
a=>a_2,
b=>"1101011100",
X=>mulr_2_836);

mulc_3_836 : entity work.gfmul
port map(
a=>a_3,
b=>"1000100110",
X=>mulr_3_836);

mulc_4_836 : entity work.gfmul
port map(
a=>a_4,
b=>"0001010101",
X=>mulr_4_836);

mulr_1_837<=a_1;
mulc_2_837 : entity work.gfmul
port map(
a=>a_2,
b=>"1010110001",
X=>mulr_2_837);

mulc_3_837 : entity work.gfmul
port map(
a=>a_3,
b=>"0010001010",
X=>mulr_3_837);

mulc_4_837 : entity work.gfmul
port map(
a=>a_4,
b=>"1010101000",
X=>mulr_4_837);

mulr_1_838<=a_1;
mulc_2_838 : entity work.gfmul
port map(
a=>a_2,
b=>"0101101011",
X=>mulr_2_838);

mulc_3_838 : entity work.gfmul
port map(
a=>a_3,
b=>"1000101000",
X=>mulr_3_838);

mulc_4_838 : entity work.gfmul
port map(
a=>a_4,
b=>"0101101101",
X=>mulr_4_838);

mulr_1_839<=a_1;
mulc_2_839 : entity work.gfmul
port map(
a=>a_2,
b=>"1011010110",
X=>mulr_2_839);

mulc_3_839 : entity work.gfmul
port map(
a=>a_3,
b=>"0010110010",
X=>mulr_3_839);

mulc_4_839 : entity work.gfmul
port map(
a=>a_4,
b=>"1101111010",
X=>mulr_4_839);

mulr_1_840<=a_1;
mulc_2_840 : entity work.gfmul
port map(
a=>a_2,
b=>"0110100101",
X=>mulr_2_840);

mulc_3_840 : entity work.gfmul
port map(
a=>a_3,
b=>"1011001000",
X=>mulr_3_840);

mulc_4_840 : entity work.gfmul
port map(
a=>a_4,
b=>"1111100110",
X=>mulr_4_840);

mulr_1_841<=a_1;
mulc_2_841 : entity work.gfmul
port map(
a=>a_2,
b=>"1101001010",
X=>mulr_2_841);

mulc_3_841 : entity work.gfmul
port map(
a=>a_3,
b=>"1100110010",
X=>mulr_3_841);

mulc_4_841 : entity work.gfmul
port map(
a=>a_4,
b=>"1100001111",
X=>mulr_4_841);

mulr_1_842<=a_1;
mulc_2_842 : entity work.gfmul
port map(
a=>a_2,
b=>"1010011101",
X=>mulr_2_842);

mulc_3_842 : entity work.gfmul
port map(
a=>a_3,
b=>"0011010011",
X=>mulr_3_842);

mulc_4_842 : entity work.gfmul
port map(
a=>a_4,
b=>"0001001110",
X=>mulr_4_842);

mulr_1_843<=a_1;
mulc_2_843 : entity work.gfmul
port map(
a=>a_2,
b=>"0100110011",
X=>mulr_2_843);

mulc_3_843 : entity work.gfmul
port map(
a=>a_3,
b=>"1101001100",
X=>mulr_3_843);

mulc_4_843 : entity work.gfmul
port map(
a=>a_4,
b=>"1001110000",
X=>mulr_4_843);

mulr_1_844<=a_1;
mulc_2_844 : entity work.gfmul
port map(
a=>a_2,
b=>"1001100110",
X=>mulr_2_844);

mulc_3_844 : entity work.gfmul
port map(
a=>a_3,
b=>"0100101011",
X=>mulr_3_844);

mulc_4_844 : entity work.gfmul
port map(
a=>a_4,
b=>"1110100100",
X=>mulr_4_844);

mulr_1_845<=a_1;
mulc_2_845 : entity work.gfmul
port map(
a=>a_2,
b=>"0011000101",
X=>mulr_2_845);

mulc_3_845 : entity work.gfmul
port map(
a=>a_3,
b=>"0010100101",
X=>mulr_3_845);

mulc_4_845 : entity work.gfmul
port map(
a=>a_4,
b=>"0100011111",
X=>mulr_4_845);

mulr_1_846<=a_1;
mulc_2_846 : entity work.gfmul
port map(
a=>a_2,
b=>"0110001010",
X=>mulr_2_846);

mulc_3_846 : entity work.gfmul
port map(
a=>a_3,
b=>"1010010100",
X=>mulr_3_846);

mulc_4_846 : entity work.gfmul
port map(
a=>a_4,
b=>"0011101010",
X=>mulr_4_846);

mulr_1_847<=a_1;
mulc_2_847 : entity work.gfmul
port map(
a=>a_2,
b=>"1100010100",
X=>mulr_2_847);

mulc_3_847 : entity work.gfmul
port map(
a=>a_3,
b=>"1001000010",
X=>mulr_3_847);

mulc_4_847 : entity work.gfmul
port map(
a=>a_4,
b=>"1101011001",
X=>mulr_4_847);

mulr_1_848<=a_1;
mulc_2_848 : entity work.gfmul
port map(
a=>a_2,
b=>"1000100001",
X=>mulr_2_848);

mulc_3_848 : entity work.gfmul
port map(
a=>a_3,
b=>"0100011010",
X=>mulr_3_848);

mulc_4_848 : entity work.gfmul
port map(
a=>a_4,
b=>"1011111110",
X=>mulr_4_848);

mulr_1_849<=a_1;
mulc_2_849 : entity work.gfmul
port map(
a=>a_2,
b=>"0001001011",
X=>mulr_2_849);

mulc_3_849 : entity work.gfmul
port map(
a=>a_3,
b=>"0001100001",
X=>mulr_3_849);

mulc_4_849 : entity work.gfmul
port map(
a=>a_4,
b=>"1111011101",
X=>mulr_4_849);

mulr_1_850<=a_1;
mulc_2_850 : entity work.gfmul
port map(
a=>a_2,
b=>"0010010110",
X=>mulr_2_850);

mulc_3_850 : entity work.gfmul
port map(
a=>a_3,
b=>"0110000100",
X=>mulr_3_850);

mulc_4_850 : entity work.gfmul
port map(
a=>a_4,
b=>"1011010111",
X=>mulr_4_850);

mulr_1_851<=a_1;
mulc_2_851 : entity work.gfmul
port map(
a=>a_2,
b=>"0100101100",
X=>mulr_2_851);

mulc_3_851 : entity work.gfmul
port map(
a=>a_3,
b=>"1000011001",
X=>mulr_3_851);

mulc_4_851 : entity work.gfmul
port map(
a=>a_4,
b=>"1010010101",
X=>mulr_4_851);

mulr_1_852<=a_1;
mulc_2_852 : entity work.gfmul
port map(
a=>a_2,
b=>"1001011000",
X=>mulr_2_852);

mulc_3_852 : entity work.gfmul
port map(
a=>a_3,
b=>"0001110110",
X=>mulr_3_852);

mulc_4_852 : entity work.gfmul
port map(
a=>a_4,
b=>"0010000101",
X=>mulr_4_852);

mulr_1_853<=a_1;
mulc_2_853 : entity work.gfmul
port map(
a=>a_2,
b=>"0010111001",
X=>mulr_2_853);

mulc_3_853 : entity work.gfmul
port map(
a=>a_3,
b=>"0111011000",
X=>mulr_3_853);

mulc_4_853 : entity work.gfmul
port map(
a=>a_4,
b=>"0000100001",
X=>mulr_4_853);

mulr_1_854<=a_1;
mulc_2_854 : entity work.gfmul
port map(
a=>a_2,
b=>"0101110010",
X=>mulr_2_854);

mulc_3_854 : entity work.gfmul
port map(
a=>a_3,
b=>"1101101001",
X=>mulr_3_854);

mulc_4_854 : entity work.gfmul
port map(
a=>a_4,
b=>"0100001000",
X=>mulr_4_854);

mulr_1_855<=a_1;
mulc_2_855 : entity work.gfmul
port map(
a=>a_2,
b=>"1011100100",
X=>mulr_2_855);

mulc_3_855 : entity work.gfmul
port map(
a=>a_3,
b=>"0110111111",
X=>mulr_3_855);

mulc_4_855 : entity work.gfmul
port map(
a=>a_4,
b=>"0001010010",
X=>mulr_4_855);

mulr_1_856<=a_1;
mulc_2_856 : entity work.gfmul
port map(
a=>a_2,
b=>"0111000001",
X=>mulr_2_856);

mulc_3_856 : entity work.gfmul
port map(
a=>a_3,
b=>"1011110101",
X=>mulr_3_856);

mulc_4_856 : entity work.gfmul
port map(
a=>a_4,
b=>"1010010000",
X=>mulr_4_856);

mulr_1_857<=a_1;
mulc_2_857 : entity work.gfmul
port map(
a=>a_2,
b=>"1110000010",
X=>mulr_2_857);

mulc_3_857 : entity work.gfmul
port map(
a=>a_3,
b=>"1111000110",
X=>mulr_3_857);

mulc_4_857 : entity work.gfmul
port map(
a=>a_4,
b=>"0010101101",
X=>mulr_4_857);

mulr_1_858<=a_1;
mulc_2_858 : entity work.gfmul
port map(
a=>a_2,
b=>"1100001101",
X=>mulr_2_858);

mulc_3_858 : entity work.gfmul
port map(
a=>a_3,
b=>"1100000011",
X=>mulr_3_858);

mulc_4_858 : entity work.gfmul
port map(
a=>a_4,
b=>"0101100001",
X=>mulr_4_858);

mulr_1_859<=a_1;
mulc_2_859 : entity work.gfmul
port map(
a=>a_2,
b=>"1000010011",
X=>mulr_2_859);

mulc_3_859 : entity work.gfmul
port map(
a=>a_3,
b=>"0000010111",
X=>mulr_3_859);

mulc_4_859 : entity work.gfmul
port map(
a=>a_4,
b=>"1100011010",
X=>mulr_4_859);

mulr_1_860<=a_1;
mulc_2_860 : entity work.gfmul
port map(
a=>a_2,
b=>"0000101111",
X=>mulr_2_860);

mulc_3_860 : entity work.gfmul
port map(
a=>a_3,
b=>"0001011100",
X=>mulr_3_860);

mulc_4_860 : entity work.gfmul
port map(
a=>a_4,
b=>"0011100110",
X=>mulr_4_860);

mulr_1_861<=a_1;
mulc_2_861 : entity work.gfmul
port map(
a=>a_2,
b=>"0001011110",
X=>mulr_2_861);

mulc_3_861 : entity work.gfmul
port map(
a=>a_3,
b=>"0101110000",
X=>mulr_3_861);

mulc_4_861 : entity work.gfmul
port map(
a=>a_4,
b=>"1100111001",
X=>mulr_4_861);

mulr_1_862<=a_1;
mulc_2_862 : entity work.gfmul
port map(
a=>a_2,
b=>"0010111100",
X=>mulr_2_862);

mulc_3_862 : entity work.gfmul
port map(
a=>a_3,
b=>"0111001001",
X=>mulr_3_862);

mulc_4_862 : entity work.gfmul
port map(
a=>a_4,
b=>"0111111110",
X=>mulr_4_862);

mulr_1_863<=a_1;
mulc_2_863 : entity work.gfmul
port map(
a=>a_2,
b=>"0101111000",
X=>mulr_2_863);

mulc_3_863 : entity work.gfmul
port map(
a=>a_3,
b=>"1100101101",
X=>mulr_3_863);

mulc_4_863 : entity work.gfmul
port map(
a=>a_4,
b=>"1111101011",
X=>mulr_4_863);

mulr_1_864<=a_1;
mulc_2_864 : entity work.gfmul
port map(
a=>a_2,
b=>"1011110000",
X=>mulr_2_864);

mulc_3_864 : entity work.gfmul
port map(
a=>a_3,
b=>"0010101111",
X=>mulr_3_864);

mulc_4_864 : entity work.gfmul
port map(
a=>a_4,
b=>"1101100111",
X=>mulr_4_864);

mulr_1_865<=a_1;
mulc_2_865 : entity work.gfmul
port map(
a=>a_2,
b=>"0111101001",
X=>mulr_2_865);

mulc_3_865 : entity work.gfmul
port map(
a=>a_3,
b=>"1010111100",
X=>mulr_3_865);

mulc_4_865 : entity work.gfmul
port map(
a=>a_4,
b=>"1100001110",
X=>mulr_4_865);

mulr_1_866<=a_1;
mulc_2_866 : entity work.gfmul
port map(
a=>a_2,
b=>"1111010010",
X=>mulr_2_866);

mulc_3_866 : entity work.gfmul
port map(
a=>a_3,
b=>"1011100010",
X=>mulr_3_866);

mulc_4_866 : entity work.gfmul
port map(
a=>a_4,
b=>"0001000110",
X=>mulr_4_866);

mulr_1_867<=a_1;
mulc_2_867 : entity work.gfmul
port map(
a=>a_2,
b=>"1110101101",
X=>mulr_2_867);

mulc_3_867 : entity work.gfmul
port map(
a=>a_3,
b=>"1110011010",
X=>mulr_3_867);

mulc_4_867 : entity work.gfmul
port map(
a=>a_4,
b=>"1000110000",
X=>mulr_4_867);

mulr_1_868<=a_1;
mulc_2_868 : entity work.gfmul
port map(
a=>a_2,
b=>"1101010011",
X=>mulr_2_868);

mulc_3_868 : entity work.gfmul
port map(
a=>a_3,
b=>"1001110011",
X=>mulr_3_868);

mulc_4_868 : entity work.gfmul
port map(
a=>a_4,
b=>"0110100100",
X=>mulr_4_868);

mulr_1_869<=a_1;
mulc_2_869 : entity work.gfmul
port map(
a=>a_2,
b=>"1010101111",
X=>mulr_2_869);

mulc_3_869 : entity work.gfmul
port map(
a=>a_3,
b=>"0111011110",
X=>mulr_3_869);

mulc_4_869 : entity work.gfmul
port map(
a=>a_4,
b=>"0100111011",
X=>mulr_4_869);

mulr_1_870<=a_1;
mulc_2_870 : entity work.gfmul
port map(
a=>a_2,
b=>"0101010111",
X=>mulr_2_870);

mulc_3_870 : entity work.gfmul
port map(
a=>a_3,
b=>"1101110001",
X=>mulr_3_870);

mulc_4_870 : entity work.gfmul
port map(
a=>a_4,
b=>"0111001010",
X=>mulr_4_870);

mulr_1_871<=a_1;
mulc_2_871 : entity work.gfmul
port map(
a=>a_2,
b=>"1010101110",
X=>mulr_2_871);

mulc_3_871 : entity work.gfmul
port map(
a=>a_3,
b=>"0111011111",
X=>mulr_3_871);

mulc_4_871 : entity work.gfmul
port map(
a=>a_4,
b=>"1001001011",
X=>mulr_4_871);

mulr_1_872<=a_1;
mulc_2_872 : entity work.gfmul
port map(
a=>a_2,
b=>"0101010101",
X=>mulr_2_872);

mulc_3_872 : entity work.gfmul
port map(
a=>a_3,
b=>"1101110101",
X=>mulr_3_872);

mulc_4_872 : entity work.gfmul
port map(
a=>a_4,
b=>"1001111100",
X=>mulr_4_872);

mulr_1_873<=a_1;
mulc_2_873 : entity work.gfmul
port map(
a=>a_2,
b=>"1010101010",
X=>mulr_2_873);

mulc_3_873 : entity work.gfmul
port map(
a=>a_3,
b=>"0111001111",
X=>mulr_3_873);

mulc_4_873 : entity work.gfmul
port map(
a=>a_4,
b=>"1111000100",
X=>mulr_4_873);

mulr_1_874<=a_1;
mulc_2_874 : entity work.gfmul
port map(
a=>a_2,
b=>"0101011101",
X=>mulr_2_874);

mulc_3_874 : entity work.gfmul
port map(
a=>a_3,
b=>"1100110101",
X=>mulr_3_874);

mulc_4_874 : entity work.gfmul
port map(
a=>a_4,
b=>"1000011111",
X=>mulr_4_874);

mulr_1_875<=a_1;
mulc_2_875 : entity work.gfmul
port map(
a=>a_2,
b=>"1010111010",
X=>mulr_2_875);

mulc_3_875 : entity work.gfmul
port map(
a=>a_3,
b=>"0011001111",
X=>mulr_3_875);

mulc_4_875 : entity work.gfmul
port map(
a=>a_4,
b=>"0011011100",
X=>mulr_4_875);

mulr_1_876<=a_1;
mulc_2_876 : entity work.gfmul
port map(
a=>a_2,
b=>"0101111101",
X=>mulr_2_876);

mulc_3_876 : entity work.gfmul
port map(
a=>a_3,
b=>"1100111100",
X=>mulr_3_876);

mulc_4_876 : entity work.gfmul
port map(
a=>a_4,
b=>"1011101001",
X=>mulr_4_876);

mulr_1_877<=a_1;
mulc_2_877 : entity work.gfmul
port map(
a=>a_2,
b=>"1011111010",
X=>mulr_2_877);

mulc_3_877 : entity work.gfmul
port map(
a=>a_3,
b=>"0011101011",
X=>mulr_3_877);

mulc_4_877 : entity work.gfmul
port map(
a=>a_4,
b=>"1101100101",
X=>mulr_4_877);

mulr_1_878<=a_1;
mulc_2_878 : entity work.gfmul
port map(
a=>a_2,
b=>"0111111101",
X=>mulr_2_878);

mulc_3_878 : entity work.gfmul
port map(
a=>a_3,
b=>"1110101100",
X=>mulr_3_878);

mulc_4_878 : entity work.gfmul
port map(
a=>a_4,
b=>"1100011110",
X=>mulr_4_878);

mulr_1_879<=a_1;
mulc_2_879 : entity work.gfmul
port map(
a=>a_2,
b=>"1111111010",
X=>mulr_2_879);

mulc_3_879 : entity work.gfmul
port map(
a=>a_3,
b=>"1010101011",
X=>mulr_3_879);

mulc_4_879 : entity work.gfmul
port map(
a=>a_4,
b=>"0011000110",
X=>mulr_4_879);

mulr_1_880<=a_1;
mulc_2_880 : entity work.gfmul
port map(
a=>a_2,
b=>"1111111101",
X=>mulr_2_880);

mulc_3_880 : entity work.gfmul
port map(
a=>a_3,
b=>"1010111110",
X=>mulr_3_880);

mulc_4_880 : entity work.gfmul
port map(
a=>a_4,
b=>"1000111001",
X=>mulr_4_880);

mulr_1_881<=a_1;
mulc_2_881 : entity work.gfmul
port map(
a=>a_2,
b=>"1111110011",
X=>mulr_2_881);

mulc_3_881 : entity work.gfmul
port map(
a=>a_3,
b=>"1011101010",
X=>mulr_3_881);

mulc_4_881 : entity work.gfmul
port map(
a=>a_4,
b=>"0111101100",
X=>mulr_4_881);

mulr_1_882<=a_1;
mulc_2_882 : entity work.gfmul
port map(
a=>a_2,
b=>"1111101111",
X=>mulr_2_882);

mulc_3_882 : entity work.gfmul
port map(
a=>a_3,
b=>"1110111010",
X=>mulr_3_882);

mulc_4_882 : entity work.gfmul
port map(
a=>a_4,
b=>"1101111011",
X=>mulr_4_882);

mulr_1_883<=a_1;
mulc_2_883 : entity work.gfmul
port map(
a=>a_2,
b=>"1111010111",
X=>mulr_2_883);

mulc_3_883 : entity work.gfmul
port map(
a=>a_3,
b=>"1011110011",
X=>mulr_3_883);

mulc_4_883 : entity work.gfmul
port map(
a=>a_4,
b=>"1111101110",
X=>mulr_4_883);

mulr_1_884<=a_1;
mulc_2_884 : entity work.gfmul
port map(
a=>a_2,
b=>"1110100111",
X=>mulr_2_884);

mulc_3_884 : entity work.gfmul
port map(
a=>a_3,
b=>"1111011110",
X=>mulr_3_884);

mulc_4_884 : entity work.gfmul
port map(
a=>a_4,
b=>"1101001111",
X=>mulr_4_884);

mulr_1_885<=a_1;
mulc_2_885 : entity work.gfmul
port map(
a=>a_2,
b=>"1101000111",
X=>mulr_2_885);

mulc_3_885 : entity work.gfmul
port map(
a=>a_3,
b=>"1101100011",
X=>mulr_3_885);

mulc_4_885 : entity work.gfmul
port map(
a=>a_4,
b=>"1001001110",
X=>mulr_4_885);

mulr_1_886<=a_1;
mulc_2_886 : entity work.gfmul
port map(
a=>a_2,
b=>"1010000111",
X=>mulr_2_886);

mulc_3_886 : entity work.gfmul
port map(
a=>a_3,
b=>"0110010111",
X=>mulr_3_886);

mulc_4_886 : entity work.gfmul
port map(
a=>a_4,
b=>"1001010100",
X=>mulr_4_886);

mulr_1_887<=a_1;
mulc_2_887 : entity work.gfmul
port map(
a=>a_2,
b=>"0100000111",
X=>mulr_2_887);

mulc_3_887 : entity work.gfmul
port map(
a=>a_3,
b=>"1001010101",
X=>mulr_3_887);

mulc_4_887 : entity work.gfmul
port map(
a=>a_4,
b=>"1010000100",
X=>mulr_4_887);

mulr_1_888<=a_1;
mulc_2_888 : entity work.gfmul
port map(
a=>a_2,
b=>"1000001110",
X=>mulr_2_888);

mulc_3_888 : entity work.gfmul
port map(
a=>a_3,
b=>"0101000110",
X=>mulr_3_888);

mulc_4_888 : entity work.gfmul
port map(
a=>a_4,
b=>"0000001101",
X=>mulr_4_888);

mulr_1_889<=a_1;
mulc_2_889 : entity work.gfmul
port map(
a=>a_2,
b=>"0000010101",
X=>mulr_2_889);

mulc_3_889 : entity work.gfmul
port map(
a=>a_3,
b=>"0100010001",
X=>mulr_3_889);

mulc_4_889 : entity work.gfmul
port map(
a=>a_4,
b=>"0001101000",
X=>mulr_4_889);

mulr_1_890<=a_1;
mulc_2_890 : entity work.gfmul
port map(
a=>a_2,
b=>"0000101010",
X=>mulr_2_890);

mulc_3_890 : entity work.gfmul
port map(
a=>a_3,
b=>"0001001101",
X=>mulr_3_890);

mulc_4_890 : entity work.gfmul
port map(
a=>a_4,
b=>"1101000000",
X=>mulr_4_890);

mulr_1_891<=a_1;
mulc_2_891 : entity work.gfmul
port map(
a=>a_2,
b=>"0001010100",
X=>mulr_2_891);

mulc_3_891 : entity work.gfmul
port map(
a=>a_3,
b=>"0100110100",
X=>mulr_3_891);

mulc_4_891 : entity work.gfmul
port map(
a=>a_4,
b=>"1000110110",
X=>mulr_4_891);

mulr_1_892<=a_1;
mulc_2_892 : entity work.gfmul
port map(
a=>a_2,
b=>"0010101000",
X=>mulr_2_892);

mulc_3_892 : entity work.gfmul
port map(
a=>a_3,
b=>"0011011001",
X=>mulr_3_892);

mulc_4_892 : entity work.gfmul
port map(
a=>a_4,
b=>"0110010100",
X=>mulr_4_892);

mulr_1_893<=a_1;
mulc_2_893 : entity work.gfmul
port map(
a=>a_2,
b=>"0101010000",
X=>mulr_2_893);

mulc_3_893 : entity work.gfmul
port map(
a=>a_3,
b=>"1101100100",
X=>mulr_3_893);

mulc_4_893 : entity work.gfmul
port map(
a=>a_4,
b=>"0010111011",
X=>mulr_4_893);

mulr_1_894<=a_1;
mulc_2_894 : entity work.gfmul
port map(
a=>a_2,
b=>"1010100000",
X=>mulr_2_894);

mulc_3_894 : entity work.gfmul
port map(
a=>a_3,
b=>"0110001011",
X=>mulr_3_894);

mulc_4_894 : entity work.gfmul
port map(
a=>a_4,
b=>"0111010001",
X=>mulr_4_894);

mulr_1_895<=a_1;
mulc_2_895 : entity work.gfmul
port map(
a=>a_2,
b=>"0101001001",
X=>mulr_2_895);

mulc_3_895 : entity work.gfmul
port map(
a=>a_3,
b=>"1000100101",
X=>mulr_3_895);

mulc_4_895 : entity work.gfmul
port map(
a=>a_4,
b=>"1010010011",
X=>mulr_4_895);

mulr_1_896<=a_1;
mulc_2_896 : entity work.gfmul
port map(
a=>a_2,
b=>"1010010010",
X=>mulr_2_896);

mulc_3_896 : entity work.gfmul
port map(
a=>a_3,
b=>"0010000110",
X=>mulr_3_896);

mulc_4_896 : entity work.gfmul
port map(
a=>a_4,
b=>"0010110101",
X=>mulr_4_896);

mulr_1_897<=a_1;
mulc_2_897 : entity work.gfmul
port map(
a=>a_2,
b=>"0100101101",
X=>mulr_2_897);

mulc_3_897 : entity work.gfmul
port map(
a=>a_3,
b=>"1000011000",
X=>mulr_3_897);

mulc_4_897 : entity work.gfmul
port map(
a=>a_4,
b=>"0110100001",
X=>mulr_4_897);

mulr_1_898<=a_1;
mulc_2_898 : entity work.gfmul
port map(
a=>a_2,
b=>"1001011010",
X=>mulr_2_898);

mulc_3_898 : entity work.gfmul
port map(
a=>a_3,
b=>"0001110010",
X=>mulr_3_898);

mulc_4_898 : entity work.gfmul
port map(
a=>a_4,
b=>"0100010011",
X=>mulr_4_898);

mulr_1_899<=a_1;
mulc_2_899 : entity work.gfmul
port map(
a=>a_2,
b=>"0010111101",
X=>mulr_2_899);

mulc_3_899 : entity work.gfmul
port map(
a=>a_3,
b=>"0111001000",
X=>mulr_3_899);

mulc_4_899 : entity work.gfmul
port map(
a=>a_4,
b=>"0010001010",
X=>mulr_4_899);

mulr_1_900<=a_1;
mulc_2_900 : entity work.gfmul
port map(
a=>a_2,
b=>"0101111010",
X=>mulr_2_900);

mulc_3_900 : entity work.gfmul
port map(
a=>a_3,
b=>"1100101001",
X=>mulr_3_900);

mulc_4_900 : entity work.gfmul
port map(
a=>a_4,
b=>"0001011001",
X=>mulr_4_900);

mulr_1_901<=a_1;
mulc_2_901 : entity work.gfmul
port map(
a=>a_2,
b=>"1011110100",
X=>mulr_2_901);

mulc_3_901 : entity work.gfmul
port map(
a=>a_3,
b=>"0010111111",
X=>mulr_3_901);

mulc_4_901 : entity work.gfmul
port map(
a=>a_4,
b=>"1011001000",
X=>mulr_4_901);

mulr_1_902<=a_1;
mulc_2_902 : entity work.gfmul
port map(
a=>a_2,
b=>"0111100001",
X=>mulr_2_902);

mulc_3_902 : entity work.gfmul
port map(
a=>a_3,
b=>"1011111100",
X=>mulr_3_902);

mulc_4_902 : entity work.gfmul
port map(
a=>a_4,
b=>"1001101101",
X=>mulr_4_902);

mulr_1_903<=a_1;
mulc_2_903 : entity work.gfmul
port map(
a=>a_2,
b=>"1111000010",
X=>mulr_2_903);

mulc_3_903 : entity work.gfmul
port map(
a=>a_3,
b=>"1111100010",
X=>mulr_3_903);

mulc_4_903 : entity work.gfmul
port map(
a=>a_4,
b=>"1101001100",
X=>mulr_4_903);

mulr_1_904<=a_1;
mulc_2_904 : entity work.gfmul
port map(
a=>a_2,
b=>"1110001101",
X=>mulr_2_904);

mulc_3_904 : entity work.gfmul
port map(
a=>a_3,
b=>"1110010011",
X=>mulr_3_904);

mulc_4_904 : entity work.gfmul
port map(
a=>a_4,
b=>"1001010110",
X=>mulr_4_904);

mulr_1_905<=a_1;
mulc_2_905 : entity work.gfmul
port map(
a=>a_2,
b=>"1100010011",
X=>mulr_2_905);

mulc_3_905 : entity work.gfmul
port map(
a=>a_3,
b=>"1001010111",
X=>mulr_3_905);

mulc_4_905 : entity work.gfmul
port map(
a=>a_4,
b=>"1010010100",
X=>mulr_4_905);

mulr_1_906<=a_1;
mulc_2_906 : entity work.gfmul
port map(
a=>a_2,
b=>"1000101111",
X=>mulr_2_906);

mulc_3_906 : entity work.gfmul
port map(
a=>a_3,
b=>"0101001110",
X=>mulr_3_906);

mulc_4_906 : entity work.gfmul
port map(
a=>a_4,
b=>"0010001101",
X=>mulr_4_906);

mulr_1_907<=a_1;
mulc_2_907 : entity work.gfmul
port map(
a=>a_2,
b=>"0001010111",
X=>mulr_2_907);

mulc_3_907 : entity work.gfmul
port map(
a=>a_3,
b=>"0100110001",
X=>mulr_3_907);

mulc_4_907 : entity work.gfmul
port map(
a=>a_4,
b=>"0001100001",
X=>mulr_4_907);

mulr_1_908<=a_1;
mulc_2_908 : entity work.gfmul
port map(
a=>a_2,
b=>"0010101110",
X=>mulr_2_908);

mulc_3_908 : entity work.gfmul
port map(
a=>a_3,
b=>"0011001101",
X=>mulr_3_908);

mulc_4_908 : entity work.gfmul
port map(
a=>a_4,
b=>"1100001000",
X=>mulr_4_908);

mulr_1_909<=a_1;
mulc_2_909 : entity work.gfmul
port map(
a=>a_2,
b=>"0101011100",
X=>mulr_2_909);

mulc_3_909 : entity work.gfmul
port map(
a=>a_3,
b=>"1100110100",
X=>mulr_3_909);

mulc_4_909 : entity work.gfmul
port map(
a=>a_4,
b=>"0001110110",
X=>mulr_4_909);

mulr_1_910<=a_1;
mulc_2_910 : entity work.gfmul
port map(
a=>a_2,
b=>"1010111000",
X=>mulr_2_910);

mulc_3_910 : entity work.gfmul
port map(
a=>a_3,
b=>"0011001011",
X=>mulr_3_910);

mulc_4_910 : entity work.gfmul
port map(
a=>a_4,
b=>"1110110000",
X=>mulr_4_910);

mulr_1_911<=a_1;
mulc_2_911 : entity work.gfmul
port map(
a=>a_2,
b=>"0101111001",
X=>mulr_2_911);

mulc_3_911 : entity work.gfmul
port map(
a=>a_3,
b=>"1100101100",
X=>mulr_3_911);

mulc_4_911 : entity work.gfmul
port map(
a=>a_4,
b=>"0110111111",
X=>mulr_4_911);

mulr_1_912<=a_1;
mulc_2_912 : entity work.gfmul
port map(
a=>a_2,
b=>"1011110010",
X=>mulr_2_912);

mulc_3_912 : entity work.gfmul
port map(
a=>a_3,
b=>"0010101011",
X=>mulr_3_912);

mulc_4_912 : entity work.gfmul
port map(
a=>a_4,
b=>"0111100011",
X=>mulr_4_912);

mulr_1_913<=a_1;
mulc_2_913 : entity work.gfmul
port map(
a=>a_2,
b=>"0111101101",
X=>mulr_2_913);

mulc_3_913 : entity work.gfmul
port map(
a=>a_3,
b=>"1010101100",
X=>mulr_3_913);

mulc_4_913 : entity work.gfmul
port map(
a=>a_4,
b=>"1100000011",
X=>mulr_4_913);

mulr_1_914<=a_1;
mulc_2_914 : entity work.gfmul
port map(
a=>a_2,
b=>"1111011010",
X=>mulr_2_914);

mulc_3_914 : entity work.gfmul
port map(
a=>a_3,
b=>"1010100010",
X=>mulr_3_914);

mulc_4_914 : entity work.gfmul
port map(
a=>a_4,
b=>"0000101110",
X=>mulr_4_914);

mulr_1_915<=a_1;
mulc_2_915 : entity work.gfmul
port map(
a=>a_2,
b=>"1110111101",
X=>mulr_2_915);

mulc_3_915 : entity work.gfmul
port map(
a=>a_3,
b=>"1010011010",
X=>mulr_3_915);

mulc_4_915 : entity work.gfmul
port map(
a=>a_4,
b=>"0101110000",
X=>mulr_4_915);

mulr_1_916<=a_1;
mulc_2_916 : entity work.gfmul
port map(
a=>a_2,
b=>"1101110011",
X=>mulr_2_916);

mulc_3_916 : entity work.gfmul
port map(
a=>a_3,
b=>"1001111010",
X=>mulr_3_916);

mulc_4_916 : entity work.gfmul
port map(
a=>a_4,
b=>"1110010010",
X=>mulr_4_916);

mulr_1_917<=a_1;
mulc_2_917 : entity work.gfmul
port map(
a=>a_2,
b=>"1011101111",
X=>mulr_2_917);

mulc_3_917 : entity work.gfmul
port map(
a=>a_3,
b=>"0111111010",
X=>mulr_3_917);

mulc_4_917 : entity work.gfmul
port map(
a=>a_4,
b=>"0010101111",
X=>mulr_4_917);

mulr_1_918<=a_1;
mulc_2_918 : entity work.gfmul
port map(
a=>a_2,
b=>"0111010111",
X=>mulr_2_918);

mulc_3_918 : entity work.gfmul
port map(
a=>a_3,
b=>"1111100001",
X=>mulr_3_918);

mulc_4_918 : entity work.gfmul
port map(
a=>a_4,
b=>"0101110001",
X=>mulr_4_918);

mulr_1_919<=a_1;
mulc_2_919 : entity work.gfmul
port map(
a=>a_2,
b=>"1110101110",
X=>mulr_2_919);

mulc_3_919 : entity work.gfmul
port map(
a=>a_3,
b=>"1110011111",
X=>mulr_3_919);

mulc_4_919 : entity work.gfmul
port map(
a=>a_4,
b=>"1110011010",
X=>mulr_4_919);

mulr_1_920<=a_1;
mulc_2_920 : entity work.gfmul
port map(
a=>a_2,
b=>"1101010101",
X=>mulr_2_920);

mulc_3_920 : entity work.gfmul
port map(
a=>a_3,
b=>"1001100111",
X=>mulr_3_920);

mulc_4_920 : entity work.gfmul
port map(
a=>a_4,
b=>"0011101111",
X=>mulr_4_920);

mulr_1_921<=a_1;
mulc_2_921 : entity work.gfmul
port map(
a=>a_2,
b=>"1010100011",
X=>mulr_2_921);

mulc_3_921 : entity work.gfmul
port map(
a=>a_3,
b=>"0110001110",
X=>mulr_3_921);

mulc_4_921 : entity work.gfmul
port map(
a=>a_4,
b=>"1101110001",
X=>mulr_4_921);

mulr_1_922<=a_1;
mulc_2_922 : entity work.gfmul
port map(
a=>a_2,
b=>"0101001111",
X=>mulr_2_922);

mulc_3_922 : entity work.gfmul
port map(
a=>a_3,
b=>"1000110001",
X=>mulr_3_922);

mulc_4_922 : entity work.gfmul
port map(
a=>a_4,
b=>"1110111110",
X=>mulr_4_922);

mulr_1_923<=a_1;
mulc_2_923 : entity work.gfmul
port map(
a=>a_2,
b=>"1010011110",
X=>mulr_2_923);

mulc_3_923 : entity work.gfmul
port map(
a=>a_3,
b=>"0011010110",
X=>mulr_3_923);

mulc_4_923 : entity work.gfmul
port map(
a=>a_4,
b=>"0111001111",
X=>mulr_4_923);

mulr_1_924<=a_1;
mulc_2_924 : entity work.gfmul
port map(
a=>a_2,
b=>"0100110101",
X=>mulr_2_924);

mulc_3_924 : entity work.gfmul
port map(
a=>a_3,
b=>"1101011000",
X=>mulr_3_924);

mulc_4_924 : entity work.gfmul
port map(
a=>a_4,
b=>"1001100011",
X=>mulr_4_924);

mulr_1_925<=a_1;
mulc_2_925 : entity work.gfmul
port map(
a=>a_2,
b=>"1001101010",
X=>mulr_2_925);

mulc_3_925 : entity work.gfmul
port map(
a=>a_3,
b=>"0101111011",
X=>mulr_3_925);

mulc_4_925 : entity work.gfmul
port map(
a=>a_4,
b=>"1100111100",
X=>mulr_4_925);

mulr_1_926<=a_1;
mulc_2_926 : entity work.gfmul
port map(
a=>a_2,
b=>"0011011101",
X=>mulr_2_926);

mulc_3_926 : entity work.gfmul
port map(
a=>a_3,
b=>"0111100101",
X=>mulr_3_926);

mulc_4_926 : entity work.gfmul
port map(
a=>a_4,
b=>"0111010110",
X=>mulr_4_926);

mulr_1_927<=a_1;
mulc_2_927 : entity work.gfmul
port map(
a=>a_2,
b=>"0110111010",
X=>mulr_2_927);

mulc_3_927 : entity work.gfmul
port map(
a=>a_3,
b=>"1110011101",
X=>mulr_3_927);

mulc_4_927 : entity work.gfmul
port map(
a=>a_4,
b=>"1010101011",
X=>mulr_4_927);

mulr_1_928<=a_1;
mulc_2_928 : entity work.gfmul
port map(
a=>a_2,
b=>"1101110100",
X=>mulr_2_928);

mulc_3_928 : entity work.gfmul
port map(
a=>a_3,
b=>"1001101111",
X=>mulr_3_928);

mulc_4_928 : entity work.gfmul
port map(
a=>a_4,
b=>"0101110101",
X=>mulr_4_928);

mulr_1_929<=a_1;
mulc_2_929 : entity work.gfmul
port map(
a=>a_2,
b=>"1011100001",
X=>mulr_2_929);

mulc_3_929 : entity work.gfmul
port map(
a=>a_3,
b=>"0110101110",
X=>mulr_3_929);

mulc_4_929 : entity work.gfmul
port map(
a=>a_4,
b=>"1110111010",
X=>mulr_4_929);

mulr_1_930<=a_1;
mulc_2_930 : entity work.gfmul
port map(
a=>a_2,
b=>"0111001011",
X=>mulr_2_930);

mulc_3_930 : entity work.gfmul
port map(
a=>a_3,
b=>"1010110001",
X=>mulr_3_930);

mulc_4_930 : entity work.gfmul
port map(
a=>a_4,
b=>"0111101111",
X=>mulr_4_930);

mulr_1_931<=a_1;
mulc_2_931 : entity work.gfmul
port map(
a=>a_2,
b=>"1110010110",
X=>mulr_2_931);

mulc_3_931 : entity work.gfmul
port map(
a=>a_3,
b=>"1011010110",
X=>mulr_3_931);

mulc_4_931 : entity work.gfmul
port map(
a=>a_4,
b=>"1101100011",
X=>mulr_4_931);

mulr_1_932<=a_1;
mulc_2_932 : entity work.gfmul
port map(
a=>a_2,
b=>"1100100101",
X=>mulr_2_932);

mulc_3_932 : entity work.gfmul
port map(
a=>a_3,
b=>"1101001010",
X=>mulr_3_932);

mulc_4_932 : entity work.gfmul
port map(
a=>a_4,
b=>"1100101110",
X=>mulr_4_932);

mulr_1_933<=a_1;
mulc_2_933 : entity work.gfmul
port map(
a=>a_2,
b=>"1001000011",
X=>mulr_2_933);

mulc_3_933 : entity work.gfmul
port map(
a=>a_3,
b=>"0100110011",
X=>mulr_3_933);

mulc_4_933 : entity work.gfmul
port map(
a=>a_4,
b=>"0101000110",
X=>mulr_4_933);

mulr_1_934<=a_1;
mulc_2_934 : entity work.gfmul
port map(
a=>a_2,
b=>"0010001111",
X=>mulr_2_934);

mulc_3_934 : entity work.gfmul
port map(
a=>a_3,
b=>"0011000101",
X=>mulr_3_934);

mulc_4_934 : entity work.gfmul
port map(
a=>a_4,
b=>"1000100010",
X=>mulr_4_934);

mulr_1_935<=a_1;
mulc_2_935 : entity work.gfmul
port map(
a=>a_2,
b=>"0100011110",
X=>mulr_2_935);

mulc_3_935 : entity work.gfmul
port map(
a=>a_3,
b=>"1100010100",
X=>mulr_3_935);

mulc_4_935 : entity work.gfmul
port map(
a=>a_4,
b=>"0100110100",
X=>mulr_4_935);

mulr_1_936<=a_1;
mulc_2_936 : entity work.gfmul
port map(
a=>a_2,
b=>"1000111100",
X=>mulr_2_936);

mulc_3_936 : entity work.gfmul
port map(
a=>a_3,
b=>"0001001011",
X=>mulr_3_936);

mulc_4_936 : entity work.gfmul
port map(
a=>a_4,
b=>"0110110010",
X=>mulr_4_936);

mulr_1_937<=a_1;
mulc_2_937 : entity work.gfmul
port map(
a=>a_2,
b=>"0001110001",
X=>mulr_2_937);

mulc_3_937 : entity work.gfmul
port map(
a=>a_3,
b=>"0100101100",
X=>mulr_3_937);

mulc_4_937 : entity work.gfmul
port map(
a=>a_4,
b=>"0110001011",
X=>mulr_4_937);

mulr_1_938<=a_1;
mulc_2_938 : entity work.gfmul
port map(
a=>a_2,
b=>"0011100010",
X=>mulr_2_938);

mulc_3_938 : entity work.gfmul
port map(
a=>a_3,
b=>"0010111001",
X=>mulr_3_938);

mulc_4_938 : entity work.gfmul
port map(
a=>a_4,
b=>"0001000011",
X=>mulr_4_938);

mulr_1_939<=a_1;
mulc_2_939 : entity work.gfmul
port map(
a=>a_2,
b=>"0111000100",
X=>mulr_2_939);

mulc_3_939 : entity work.gfmul
port map(
a=>a_3,
b=>"1011100100",
X=>mulr_3_939);

mulc_4_939 : entity work.gfmul
port map(
a=>a_4,
b=>"1000011000",
X=>mulr_4_939);

mulr_1_940<=a_1;
mulc_2_940 : entity work.gfmul
port map(
a=>a_2,
b=>"1110001000",
X=>mulr_2_940);

mulc_3_940 : entity work.gfmul
port map(
a=>a_3,
b=>"1110000010",
X=>mulr_3_940);

mulc_4_940 : entity work.gfmul
port map(
a=>a_4,
b=>"0011100100",
X=>mulr_4_940);

mulr_1_941<=a_1;
mulc_2_941 : entity work.gfmul
port map(
a=>a_2,
b=>"1100011001",
X=>mulr_2_941);

mulc_3_941 : entity work.gfmul
port map(
a=>a_3,
b=>"1000010011",
X=>mulr_3_941);

mulc_4_941 : entity work.gfmul
port map(
a=>a_4,
b=>"1100101001",
X=>mulr_4_941);

mulr_1_942<=a_1;
mulc_2_942 : entity work.gfmul
port map(
a=>a_2,
b=>"1000111011",
X=>mulr_2_942);

mulc_3_942 : entity work.gfmul
port map(
a=>a_3,
b=>"0001011110",
X=>mulr_3_942);

mulc_4_942 : entity work.gfmul
port map(
a=>a_4,
b=>"0101111110",
X=>mulr_4_942);

mulr_1_943<=a_1;
mulc_2_943 : entity work.gfmul
port map(
a=>a_2,
b=>"0001111111",
X=>mulr_2_943);

mulc_3_943 : entity work.gfmul
port map(
a=>a_3,
b=>"0101111000",
X=>mulr_3_943);

mulc_4_943 : entity work.gfmul
port map(
a=>a_4,
b=>"1111100010",
X=>mulr_4_943);

mulr_1_944<=a_1;
mulc_2_944 : entity work.gfmul
port map(
a=>a_2,
b=>"0011111110",
X=>mulr_2_944);

mulc_3_944 : entity work.gfmul
port map(
a=>a_3,
b=>"0111101001",
X=>mulr_3_944);

mulc_4_944 : entity work.gfmul
port map(
a=>a_4,
b=>"1100101111",
X=>mulr_4_944);

mulr_1_945<=a_1;
mulc_2_945 : entity work.gfmul
port map(
a=>a_2,
b=>"0111111100",
X=>mulr_2_945);

mulc_3_945 : entity work.gfmul
port map(
a=>a_3,
b=>"1110101101",
X=>mulr_3_945);

mulc_4_945 : entity work.gfmul
port map(
a=>a_4,
b=>"0101001110",
X=>mulr_4_945);

mulr_1_946<=a_1;
mulc_2_946 : entity work.gfmul
port map(
a=>a_2,
b=>"1111111000",
X=>mulr_2_946);

mulc_3_946 : entity work.gfmul
port map(
a=>a_3,
b=>"1010101111",
X=>mulr_3_946);

mulc_4_946 : entity work.gfmul
port map(
a=>a_4,
b=>"1001100010",
X=>mulr_4_946);

mulr_1_947<=a_1;
mulc_2_947 : entity work.gfmul
port map(
a=>a_2,
b=>"1111111001",
X=>mulr_2_947);

mulc_3_947 : entity work.gfmul
port map(
a=>a_3,
b=>"1010101110",
X=>mulr_3_947);

mulc_4_947 : entity work.gfmul
port map(
a=>a_4,
b=>"1100110100",
X=>mulr_4_947);

mulr_1_948<=a_1;
mulc_2_948 : entity work.gfmul
port map(
a=>a_2,
b=>"1111111011",
X=>mulr_2_948);

mulc_3_948 : entity work.gfmul
port map(
a=>a_3,
b=>"1010101010",
X=>mulr_3_948);

mulc_4_948 : entity work.gfmul
port map(
a=>a_4,
b=>"0110010110",
X=>mulr_4_948);

mulr_1_949<=a_1;
mulc_2_949 : entity work.gfmul
port map(
a=>a_2,
b=>"1111111111",
X=>mulr_2_949);

mulc_3_949 : entity work.gfmul
port map(
a=>a_3,
b=>"1010111010",
X=>mulr_3_949);

mulc_4_949 : entity work.gfmul
port map(
a=>a_4,
b=>"0010101011",
X=>mulr_4_949);

mulr_1_950<=a_1;
mulc_2_950 : entity work.gfmul
port map(
a=>a_2,
b=>"1111110111",
X=>mulr_2_950);

mulc_3_950 : entity work.gfmul
port map(
a=>a_3,
b=>"1011111010",
X=>mulr_3_950);

mulc_4_950 : entity work.gfmul
port map(
a=>a_4,
b=>"0101010001",
X=>mulr_4_950);

mulr_1_951<=a_1;
mulc_2_951 : entity work.gfmul
port map(
a=>a_2,
b=>"1111100111",
X=>mulr_2_951);

mulc_3_951 : entity work.gfmul
port map(
a=>a_3,
b=>"1111111010",
X=>mulr_3_951);

mulc_4_951 : entity work.gfmul
port map(
a=>a_4,
b=>"1010011010",
X=>mulr_4_951);

mulr_1_952<=a_1;
mulc_2_952 : entity work.gfmul
port map(
a=>a_2,
b=>"1111000111",
X=>mulr_2_952);

mulc_3_952 : entity work.gfmul
port map(
a=>a_3,
b=>"1111110011",
X=>mulr_3_952);

mulc_4_952 : entity work.gfmul
port map(
a=>a_4,
b=>"0011111101",
X=>mulr_4_952);

mulr_1_953<=a_1;
mulc_2_953 : entity work.gfmul
port map(
a=>a_2,
b=>"1110000111",
X=>mulr_2_953);

mulc_3_953 : entity work.gfmul
port map(
a=>a_3,
b=>"1111010111",
X=>mulr_3_953);

mulc_4_953 : entity work.gfmul
port map(
a=>a_4,
b=>"1111100001",
X=>mulr_4_953);

mulr_1_954<=a_1;
mulc_2_954 : entity work.gfmul
port map(
a=>a_2,
b=>"1100000111",
X=>mulr_2_954);

mulc_3_954 : entity work.gfmul
port map(
a=>a_3,
b=>"1101000111",
X=>mulr_3_954);

mulc_4_954 : entity work.gfmul
port map(
a=>a_4,
b=>"1100110111",
X=>mulr_4_954);

mulr_1_955<=a_1;
mulc_2_955 : entity work.gfmul
port map(
a=>a_2,
b=>"1000000111",
X=>mulr_2_955);

mulc_3_955 : entity work.gfmul
port map(
a=>a_3,
b=>"0100000111",
X=>mulr_3_955);

mulc_4_955 : entity work.gfmul
port map(
a=>a_4,
b=>"0110001110",
X=>mulr_4_955);

mulr_1_956<=a_1;
mulc_2_956 : entity work.gfmul
port map(
a=>a_2,
b=>"0000000111",
X=>mulr_2_956);

mulc_3_956 : entity work.gfmul
port map(
a=>a_3,
b=>"0000010101",
X=>mulr_3_956);

mulc_4_956 : entity work.gfmul
port map(
a=>a_4,
b=>"0001101011",
X=>mulr_4_956);

mulr_1_957<=a_1;
mulc_2_957 : entity work.gfmul
port map(
a=>a_2,
b=>"0000001110",
X=>mulr_2_957);

mulc_3_957 : entity work.gfmul
port map(
a=>a_3,
b=>"0001010100",
X=>mulr_3_957);

mulc_4_957 : entity work.gfmul
port map(
a=>a_4,
b=>"1101011000",
X=>mulr_4_957);

mulr_1_958<=a_1;
mulc_2_958 : entity work.gfmul
port map(
a=>a_2,
b=>"0000011100",
X=>mulr_2_958);

mulc_3_958 : entity work.gfmul
port map(
a=>a_3,
b=>"0101010000",
X=>mulr_3_958);

mulc_4_958 : entity work.gfmul
port map(
a=>a_4,
b=>"1011110110",
X=>mulr_4_958);

mulr_1_959<=a_1;
mulc_2_959 : entity work.gfmul
port map(
a=>a_2,
b=>"0000111000",
X=>mulr_2_959);

mulc_3_959 : entity work.gfmul
port map(
a=>a_3,
b=>"0101001001",
X=>mulr_3_959);

mulc_4_959 : entity work.gfmul
port map(
a=>a_4,
b=>"1110011101",
X=>mulr_4_959);

mulr_1_960<=a_1;
mulc_2_960 : entity work.gfmul
port map(
a=>a_2,
b=>"0001110000",
X=>mulr_2_960);

mulc_3_960 : entity work.gfmul
port map(
a=>a_3,
b=>"0100101101",
X=>mulr_3_960);

mulc_4_960 : entity work.gfmul
port map(
a=>a_4,
b=>"0011010111",
X=>mulr_4_960);

mulr_1_961<=a_1;
mulc_2_961 : entity work.gfmul
port map(
a=>a_2,
b=>"0011100000",
X=>mulr_2_961);

mulc_3_961 : entity work.gfmul
port map(
a=>a_3,
b=>"0010111101",
X=>mulr_3_961);

mulc_4_961 : entity work.gfmul
port map(
a=>a_4,
b=>"1010110001",
X=>mulr_4_961);

mulr_1_962<=a_1;
mulc_2_962 : entity work.gfmul
port map(
a=>a_2,
b=>"0111000000",
X=>mulr_2_962);

mulc_3_962 : entity work.gfmul
port map(
a=>a_3,
b=>"1011110100",
X=>mulr_3_962);

mulc_4_962 : entity work.gfmul
port map(
a=>a_4,
b=>"0110100101",
X=>mulr_4_962);

mulr_1_963<=a_1;
mulc_2_963 : entity work.gfmul
port map(
a=>a_2,
b=>"1110000000",
X=>mulr_2_963);

mulc_3_963 : entity work.gfmul
port map(
a=>a_3,
b=>"1111000010",
X=>mulr_3_963);

mulc_4_963 : entity work.gfmul
port map(
a=>a_4,
b=>"0100110011",
X=>mulr_4_963);

mulr_1_964<=a_1;
mulc_2_964 : entity work.gfmul
port map(
a=>a_2,
b=>"1100001001",
X=>mulr_2_964);

mulc_3_964 : entity work.gfmul
port map(
a=>a_3,
b=>"1100010011",
X=>mulr_3_964);

mulc_4_964 : entity work.gfmul
port map(
a=>a_4,
b=>"0110001010",
X=>mulr_4_964);

mulr_1_965<=a_1;
mulc_2_965 : entity work.gfmul
port map(
a=>a_2,
b=>"1000011011",
X=>mulr_2_965);

mulc_3_965 : entity work.gfmul
port map(
a=>a_3,
b=>"0001010111",
X=>mulr_3_965);

mulc_4_965 : entity work.gfmul
port map(
a=>a_4,
b=>"0001001011",
X=>mulr_4_965);

mulr_1_966<=a_1;
mulc_2_966 : entity work.gfmul
port map(
a=>a_2,
b=>"0000111111",
X=>mulr_2_966);

mulc_3_966 : entity work.gfmul
port map(
a=>a_3,
b=>"0101011100",
X=>mulr_3_966);

mulc_4_966 : entity work.gfmul
port map(
a=>a_4,
b=>"1001011000",
X=>mulr_4_966);

mulr_1_967<=a_1;
mulc_2_967 : entity work.gfmul
port map(
a=>a_2,
b=>"0001111110",
X=>mulr_2_967);

mulc_3_967 : entity work.gfmul
port map(
a=>a_3,
b=>"0101111001",
X=>mulr_3_967);

mulc_4_967 : entity work.gfmul
port map(
a=>a_4,
b=>"1011100100",
X=>mulr_4_967);

mulr_1_968<=a_1;
mulc_2_968 : entity work.gfmul
port map(
a=>a_2,
b=>"0011111100",
X=>mulr_2_968);

mulc_3_968 : entity work.gfmul
port map(
a=>a_3,
b=>"0111101101",
X=>mulr_3_968);

mulc_4_968 : entity work.gfmul
port map(
a=>a_4,
b=>"1100001101",
X=>mulr_4_968);

mulr_1_969<=a_1;
mulc_2_969 : entity work.gfmul
port map(
a=>a_2,
b=>"0111111000",
X=>mulr_2_969);

mulc_3_969 : entity work.gfmul
port map(
a=>a_3,
b=>"1110111101",
X=>mulr_3_969);

mulc_4_969 : entity work.gfmul
port map(
a=>a_4,
b=>"0001011110",
X=>mulr_4_969);

mulr_1_970<=a_1;
mulc_2_970 : entity work.gfmul
port map(
a=>a_2,
b=>"1111110000",
X=>mulr_2_970);

mulc_3_970 : entity work.gfmul
port map(
a=>a_3,
b=>"1011101111",
X=>mulr_3_970);

mulc_4_970 : entity work.gfmul
port map(
a=>a_4,
b=>"1011110000",
X=>mulr_4_970);

mulr_1_971<=a_1;
mulc_2_971 : entity work.gfmul
port map(
a=>a_2,
b=>"1111101001",
X=>mulr_2_971);

mulc_3_971 : entity work.gfmul
port map(
a=>a_3,
b=>"1110101110",
X=>mulr_3_971);

mulc_4_971 : entity work.gfmul
port map(
a=>a_4,
b=>"1110101101",
X=>mulr_4_971);

mulr_1_972<=a_1;
mulc_2_972 : entity work.gfmul
port map(
a=>a_2,
b=>"1111011011",
X=>mulr_2_972);

mulc_3_972 : entity work.gfmul
port map(
a=>a_3,
b=>"1010100011",
X=>mulr_3_972);

mulc_4_972 : entity work.gfmul
port map(
a=>a_4,
b=>"0101010111",
X=>mulr_4_972);

mulr_1_973<=a_1;
mulc_2_973 : entity work.gfmul
port map(
a=>a_2,
b=>"1110111111",
X=>mulr_2_973);

mulc_3_973 : entity work.gfmul
port map(
a=>a_3,
b=>"1010011110",
X=>mulr_3_973);

mulc_4_973 : entity work.gfmul
port map(
a=>a_4,
b=>"1010101010",
X=>mulr_4_973);

mulr_1_974<=a_1;
mulc_2_974 : entity work.gfmul
port map(
a=>a_2,
b=>"1101110111",
X=>mulr_2_974);

mulc_3_974 : entity work.gfmul
port map(
a=>a_3,
b=>"1001101010",
X=>mulr_3_974);

mulc_4_974 : entity work.gfmul
port map(
a=>a_4,
b=>"0101111101",
X=>mulr_4_974);

mulr_1_975<=a_1;
mulc_2_975 : entity work.gfmul
port map(
a=>a_2,
b=>"1011100111",
X=>mulr_2_975);

mulc_3_975 : entity work.gfmul
port map(
a=>a_3,
b=>"0110111010",
X=>mulr_3_975);

mulc_4_975 : entity work.gfmul
port map(
a=>a_4,
b=>"1111111010",
X=>mulr_4_975);

mulr_1_976<=a_1;
mulc_2_976 : entity work.gfmul
port map(
a=>a_2,
b=>"0111000111",
X=>mulr_2_976);

mulc_3_976 : entity work.gfmul
port map(
a=>a_3,
b=>"1011100001",
X=>mulr_3_976);

mulc_4_976 : entity work.gfmul
port map(
a=>a_4,
b=>"1111101111",
X=>mulr_4_976);

mulr_1_977<=a_1;
mulc_2_977 : entity work.gfmul
port map(
a=>a_2,
b=>"1110001110",
X=>mulr_2_977);

mulc_3_977 : entity work.gfmul
port map(
a=>a_3,
b=>"1110010110",
X=>mulr_3_977);

mulc_4_977 : entity work.gfmul
port map(
a=>a_4,
b=>"1101000111",
X=>mulr_4_977);

mulr_1_978<=a_1;
mulc_2_978 : entity work.gfmul
port map(
a=>a_2,
b=>"1100010101",
X=>mulr_2_978);

mulc_3_978 : entity work.gfmul
port map(
a=>a_3,
b=>"1001000011",
X=>mulr_3_978);

mulc_4_978 : entity work.gfmul
port map(
a=>a_4,
b=>"1000001110",
X=>mulr_4_978);

mulr_1_979<=a_1;
mulc_2_979 : entity work.gfmul
port map(
a=>a_2,
b=>"1000100011",
X=>mulr_2_979);

mulc_3_979 : entity work.gfmul
port map(
a=>a_3,
b=>"0100011110",
X=>mulr_3_979);

mulc_4_979 : entity work.gfmul
port map(
a=>a_4,
b=>"0001010100",
X=>mulr_4_979);

mulr_1_980<=a_1;
mulc_2_980 : entity work.gfmul
port map(
a=>a_2,
b=>"0001001111",
X=>mulr_2_980);

mulc_3_980 : entity work.gfmul
port map(
a=>a_3,
b=>"0001110001",
X=>mulr_3_980);

mulc_4_980 : entity work.gfmul
port map(
a=>a_4,
b=>"1010100000",
X=>mulr_4_980);

mulr_1_981<=a_1;
mulc_2_981 : entity work.gfmul
port map(
a=>a_2,
b=>"0010011110",
X=>mulr_2_981);

mulc_3_981 : entity work.gfmul
port map(
a=>a_3,
b=>"0111000100",
X=>mulr_3_981);

mulc_4_981 : entity work.gfmul
port map(
a=>a_4,
b=>"0100101101",
X=>mulr_4_981);

mulr_1_982<=a_1;
mulc_2_982 : entity work.gfmul
port map(
a=>a_2,
b=>"0100111100",
X=>mulr_2_982);

mulc_3_982 : entity work.gfmul
port map(
a=>a_3,
b=>"1100011001",
X=>mulr_3_982);

mulc_4_982 : entity work.gfmul
port map(
a=>a_4,
b=>"0101111010",
X=>mulr_4_982);

mulr_1_983<=a_1;
mulc_2_983 : entity work.gfmul
port map(
a=>a_2,
b=>"1001111000",
X=>mulr_2_983);

mulc_3_983 : entity work.gfmul
port map(
a=>a_3,
b=>"0001111111",
X=>mulr_3_983);

mulc_4_983 : entity work.gfmul
port map(
a=>a_4,
b=>"1111000010",
X=>mulr_4_983);

mulr_1_984<=a_1;
mulc_2_984 : entity work.gfmul
port map(
a=>a_2,
b=>"0011111001",
X=>mulr_2_984);

mulc_3_984 : entity work.gfmul
port map(
a=>a_3,
b=>"0111111100",
X=>mulr_3_984);

mulc_4_984 : entity work.gfmul
port map(
a=>a_4,
b=>"1000101111",
X=>mulr_4_984);

mulr_1_985<=a_1;
mulc_2_985 : entity work.gfmul
port map(
a=>a_2,
b=>"0111110010",
X=>mulr_2_985);

mulc_3_985 : entity work.gfmul
port map(
a=>a_3,
b=>"1111111001",
X=>mulr_3_985);

mulc_4_985 : entity work.gfmul
port map(
a=>a_4,
b=>"0101011100",
X=>mulr_4_985);

mulr_1_986<=a_1;
mulc_2_986 : entity work.gfmul
port map(
a=>a_2,
b=>"1111100100",
X=>mulr_2_986);

mulc_3_986 : entity work.gfmul
port map(
a=>a_3,
b=>"1111111111",
X=>mulr_3_986);

mulc_4_986 : entity work.gfmul
port map(
a=>a_4,
b=>"1011110010",
X=>mulr_4_986);

mulr_1_987<=a_1;
mulc_2_987 : entity work.gfmul
port map(
a=>a_2,
b=>"1111000001",
X=>mulr_2_987);

mulc_3_987 : entity work.gfmul
port map(
a=>a_3,
b=>"1111100111",
X=>mulr_3_987);

mulc_4_987 : entity work.gfmul
port map(
a=>a_4,
b=>"1110111101",
X=>mulr_4_987);

mulr_1_988<=a_1;
mulc_2_988 : entity work.gfmul
port map(
a=>a_2,
b=>"1110001011",
X=>mulr_2_988);

mulc_3_988 : entity work.gfmul
port map(
a=>a_3,
b=>"1110000111",
X=>mulr_3_988);

mulc_4_988 : entity work.gfmul
port map(
a=>a_4,
b=>"0111010111",
X=>mulr_4_988);

mulr_1_989<=a_1;
mulc_2_989 : entity work.gfmul
port map(
a=>a_2,
b=>"1100011111",
X=>mulr_2_989);

mulc_3_989 : entity work.gfmul
port map(
a=>a_3,
b=>"1000000111",
X=>mulr_3_989);

mulc_4_989 : entity work.gfmul
port map(
a=>a_4,
b=>"1010100011",
X=>mulr_4_989);

mulr_1_990<=a_1;
mulc_2_990 : entity work.gfmul
port map(
a=>a_2,
b=>"1000110111",
X=>mulr_2_990);

mulc_3_990 : entity work.gfmul
port map(
a=>a_3,
b=>"0000001110",
X=>mulr_3_990);

mulc_4_990 : entity work.gfmul
port map(
a=>a_4,
b=>"0100110101",
X=>mulr_4_990);

mulr_1_991<=a_1;
mulc_2_991 : entity work.gfmul
port map(
a=>a_2,
b=>"0001100111",
X=>mulr_2_991);

mulc_3_991 : entity work.gfmul
port map(
a=>a_3,
b=>"0000111000",
X=>mulr_3_991);

mulc_4_991 : entity work.gfmul
port map(
a=>a_4,
b=>"0110111010",
X=>mulr_4_991);

mulr_1_992<=a_1;
mulc_2_992 : entity work.gfmul
port map(
a=>a_2,
b=>"0011001110",
X=>mulr_2_992);

mulc_3_992 : entity work.gfmul
port map(
a=>a_3,
b=>"0011100000",
X=>mulr_3_992);

mulc_4_992 : entity work.gfmul
port map(
a=>a_4,
b=>"0111001011",
X=>mulr_4_992);

mulr_1_993<=a_1;
mulc_2_993 : entity work.gfmul
port map(
a=>a_2,
b=>"0110011100",
X=>mulr_2_993);

mulc_3_993 : entity work.gfmul
port map(
a=>a_3,
b=>"1110000000",
X=>mulr_3_993);

mulc_4_993 : entity work.gfmul
port map(
a=>a_4,
b=>"1001000011",
X=>mulr_4_993);

mulr_1_994<=a_1;
mulc_2_994 : entity work.gfmul
port map(
a=>a_2,
b=>"1100111000",
X=>mulr_2_994);

mulc_3_994 : entity work.gfmul
port map(
a=>a_3,
b=>"1000011011",
X=>mulr_3_994);

mulc_4_994 : entity work.gfmul
port map(
a=>a_4,
b=>"1000111100",
X=>mulr_4_994);

mulr_1_995<=a_1;
mulc_2_995 : entity work.gfmul
port map(
a=>a_2,
b=>"1001111001",
X=>mulr_2_995);

mulc_3_995 : entity work.gfmul
port map(
a=>a_3,
b=>"0001111110",
X=>mulr_3_995);

mulc_4_995 : entity work.gfmul
port map(
a=>a_4,
b=>"0111000100",
X=>mulr_4_995);

mulr_1_996<=a_1;
mulc_2_996 : entity work.gfmul
port map(
a=>a_2,
b=>"0011111011",
X=>mulr_2_996);

mulc_3_996 : entity work.gfmul
port map(
a=>a_3,
b=>"0111111000",
X=>mulr_3_996);

mulc_4_996 : entity work.gfmul
port map(
a=>a_4,
b=>"1000111011",
X=>mulr_4_996);

mulr_1_997<=a_1;
mulc_2_997 : entity work.gfmul
port map(
a=>a_2,
b=>"0111110110",
X=>mulr_2_997);

mulc_3_997 : entity work.gfmul
port map(
a=>a_3,
b=>"1111101001",
X=>mulr_3_997);

mulc_4_997 : entity work.gfmul
port map(
a=>a_4,
b=>"0111111100",
X=>mulr_4_997);

mulr_1_998<=a_1;
mulc_2_998 : entity work.gfmul
port map(
a=>a_2,
b=>"1111101100",
X=>mulr_2_998);

mulc_3_998 : entity work.gfmul
port map(
a=>a_3,
b=>"1110111111",
X=>mulr_3_998);

mulc_4_998 : entity work.gfmul
port map(
a=>a_4,
b=>"1111111011",
X=>mulr_4_998);

mulr_1_999<=a_1;
mulc_2_999 : entity work.gfmul
port map(
a=>a_2,
b=>"1111010001",
X=>mulr_2_999);

mulc_3_999 : entity work.gfmul
port map(
a=>a_3,
b=>"1011100111",
X=>mulr_3_999);

mulc_4_999 : entity work.gfmul
port map(
a=>a_4,
b=>"1111100111",
X=>mulr_4_999);

mulr_1_1000<=a_1;
mulc_2_1000 : entity work.gfmul
port map(
a=>a_2,
b=>"1110101011",
X=>mulr_2_1000);

mulc_3_1000 : entity work.gfmul
port map(
a=>a_3,
b=>"1110001110",
X=>mulr_3_1000);

mulc_4_1000 : entity work.gfmul
port map(
a=>a_4,
b=>"1100000111",
X=>mulr_4_1000);

mulr_1_1001<=a_1;
mulc_2_1001 : entity work.gfmul
port map(
a=>a_2,
b=>"1101011111",
X=>mulr_2_1001);

mulc_3_1001 : entity work.gfmul
port map(
a=>a_3,
b=>"1000100011",
X=>mulr_3_1001);

mulc_4_1001 : entity work.gfmul
port map(
a=>a_4,
b=>"0000001110",
X=>mulr_4_1001);

mulr_1_1002<=a_1;
mulc_2_1002 : entity work.gfmul
port map(
a=>a_2,
b=>"1010110111",
X=>mulr_2_1002);

mulc_3_1002 : entity work.gfmul
port map(
a=>a_3,
b=>"0010011110",
X=>mulr_3_1002);

mulc_4_1002 : entity work.gfmul
port map(
a=>a_4,
b=>"0001110000",
X=>mulr_4_1002);

mulr_1_1003<=a_1;
mulc_2_1003 : entity work.gfmul
port map(
a=>a_2,
b=>"0101100111",
X=>mulr_2_1003);

mulc_3_1003 : entity work.gfmul
port map(
a=>a_3,
b=>"1001111000",
X=>mulr_3_1003);

mulc_4_1003 : entity work.gfmul
port map(
a=>a_4,
b=>"1110000000",
X=>mulr_4_1003);

mulr_1_1004<=a_1;
mulc_2_1004 : entity work.gfmul
port map(
a=>a_2,
b=>"1011001110",
X=>mulr_2_1004);

mulc_3_1004 : entity work.gfmul
port map(
a=>a_3,
b=>"0111110010",
X=>mulr_3_1004);

mulc_4_1004 : entity work.gfmul
port map(
a=>a_4,
b=>"0000111111",
X=>mulr_4_1004);

mulr_1_1005<=a_1;
mulc_2_1005 : entity work.gfmul
port map(
a=>a_2,
b=>"0110010101",
X=>mulr_2_1005);

mulc_3_1005 : entity work.gfmul
port map(
a=>a_3,
b=>"1111000001",
X=>mulr_3_1005);

mulc_4_1005 : entity work.gfmul
port map(
a=>a_4,
b=>"0111111000",
X=>mulr_4_1005);

mulr_1_1006<=a_1;
mulc_2_1006 : entity work.gfmul
port map(
a=>a_2,
b=>"1100101010",
X=>mulr_2_1006);

mulc_3_1006 : entity work.gfmul
port map(
a=>a_3,
b=>"1100011111",
X=>mulr_3_1006);

mulc_4_1006 : entity work.gfmul
port map(
a=>a_4,
b=>"1111011011",
X=>mulr_4_1006);

mulr_1_1007<=a_1;
mulc_2_1007 : entity work.gfmul
port map(
a=>a_2,
b=>"1001011101",
X=>mulr_2_1007);

mulc_3_1007 : entity work.gfmul
port map(
a=>a_3,
b=>"0001100111",
X=>mulr_3_1007);

mulc_4_1007 : entity work.gfmul
port map(
a=>a_4,
b=>"1011100111",
X=>mulr_4_1007);

mulr_1_1008<=a_1;
mulc_2_1008 : entity work.gfmul
port map(
a=>a_2,
b=>"0010110011",
X=>mulr_2_1008);

mulc_3_1008 : entity work.gfmul
port map(
a=>a_3,
b=>"0110011100",
X=>mulr_3_1008);

mulc_4_1008 : entity work.gfmul
port map(
a=>a_4,
b=>"1100010101",
X=>mulr_4_1008);

mulr_1_1009<=a_1;
mulc_2_1009 : entity work.gfmul
port map(
a=>a_2,
b=>"0101100110",
X=>mulr_2_1009);

mulc_3_1009 : entity work.gfmul
port map(
a=>a_3,
b=>"1001111001",
X=>mulr_3_1009);

mulc_4_1009 : entity work.gfmul
port map(
a=>a_4,
b=>"0010011110",
X=>mulr_4_1009);

mulr_1_1010<=a_1;
mulc_2_1010 : entity work.gfmul
port map(
a=>a_2,
b=>"1011001100",
X=>mulr_2_1010);

mulc_3_1010 : entity work.gfmul
port map(
a=>a_3,
b=>"0111110110",
X=>mulr_3_1010);

mulc_4_1010 : entity work.gfmul
port map(
a=>a_4,
b=>"0011111001",
X=>mulr_4_1010);

mulr_1_1011<=a_1;
mulc_2_1011 : entity work.gfmul
port map(
a=>a_2,
b=>"0110010001",
X=>mulr_2_1011);

mulc_3_1011 : entity work.gfmul
port map(
a=>a_3,
b=>"1111010001",
X=>mulr_3_1011);

mulc_4_1011 : entity work.gfmul
port map(
a=>a_4,
b=>"1111000001",
X=>mulr_4_1011);

mulr_1_1012<=a_1;
mulc_2_1012 : entity work.gfmul
port map(
a=>a_2,
b=>"1100100010",
X=>mulr_2_1012);

mulc_3_1012 : entity work.gfmul
port map(
a=>a_3,
b=>"1101011111",
X=>mulr_3_1012);

mulc_4_1012 : entity work.gfmul
port map(
a=>a_4,
b=>"1000110111",
X=>mulr_4_1012);

mulr_1_1013<=a_1;
mulc_2_1013 : entity work.gfmul
port map(
a=>a_2,
b=>"1001001101",
X=>mulr_2_1013);

mulc_3_1013 : entity work.gfmul
port map(
a=>a_3,
b=>"0101100111",
X=>mulr_3_1013);

mulc_4_1013 : entity work.gfmul
port map(
a=>a_4,
b=>"0110011100",
X=>mulr_4_1013);

mulr_1_1014<=a_1;
mulc_2_1014 : entity work.gfmul
port map(
a=>a_2,
b=>"0010010011",
X=>mulr_2_1014);

mulc_3_1014 : entity work.gfmul
port map(
a=>a_3,
b=>"0110010101",
X=>mulr_3_1014);

mulc_4_1014 : entity work.gfmul
port map(
a=>a_4,
b=>"0011111011",
X=>mulr_4_1014);

mulr_1_1015<=a_1;
mulc_2_1015 : entity work.gfmul
port map(
a=>a_2,
b=>"0100100110",
X=>mulr_2_1015);

mulc_3_1015 : entity work.gfmul
port map(
a=>a_3,
b=>"1001011101",
X=>mulr_3_1015);

mulc_4_1015 : entity work.gfmul
port map(
a=>a_4,
b=>"1111010001",
X=>mulr_4_1015);

mulr_1_1016<=a_1;
mulc_2_1016 : entity work.gfmul
port map(
a=>a_2,
b=>"1001001100",
X=>mulr_2_1016);

mulc_3_1016 : entity work.gfmul
port map(
a=>a_3,
b=>"0101100110",
X=>mulr_3_1016);

mulc_4_1016 : entity work.gfmul
port map(
a=>a_4,
b=>"1010110111",
X=>mulr_4_1016);

mulr_1_1017<=a_1;
mulc_2_1017 : entity work.gfmul
port map(
a=>a_2,
b=>"0010010001",
X=>mulr_2_1017);

mulc_3_1017 : entity work.gfmul
port map(
a=>a_3,
b=>"0110010001",
X=>mulr_3_1017);

mulc_4_1017 : entity work.gfmul
port map(
a=>a_4,
b=>"0110010101",
X=>mulr_4_1017);

mulr_1_1018<=a_1;
mulc_2_1018 : entity work.gfmul
port map(
a=>a_2,
b=>"0100100010",
X=>mulr_2_1018);

mulc_3_1018 : entity work.gfmul
port map(
a=>a_3,
b=>"1001001101",
X=>mulr_3_1018);

mulc_4_1018 : entity work.gfmul
port map(
a=>a_4,
b=>"0010110011",
X=>mulr_4_1018);

mulr_1_1019<=a_1;
mulc_2_1019 : entity work.gfmul
port map(
a=>a_2,
b=>"1001000100",
X=>mulr_2_1019);

mulc_3_1019 : entity work.gfmul
port map(
a=>a_3,
b=>"0100100110",
X=>mulr_3_1019);

mulc_4_1019 : entity work.gfmul
port map(
a=>a_4,
b=>"0110010001",
X=>mulr_4_1019);

mulr_1_1020<=a_1;
mulc_2_1020 : entity work.gfmul
port map(
a=>a_2,
b=>"0010000001",
X=>mulr_2_1020);

mulc_3_1020 : entity work.gfmul
port map(
a=>a_3,
b=>"0010010001",
X=>mulr_3_1020);

mulc_4_1020 : entity work.gfmul
port map(
a=>a_4,
b=>"0010010011",
X=>mulr_4_1020);

mulr_1_1021<=a_1;
mulc_2_1021 : entity work.gfmul
port map(
a=>a_2,
b=>"0100000010",
X=>mulr_2_1021);

mulc_3_1021 : entity work.gfmul
port map(
a=>a_3,
b=>"1001000100",
X=>mulr_3_1021);

mulc_4_1021 : entity work.gfmul
port map(
a=>a_4,
b=>"0010010001",
X=>mulr_4_1021);

mulr_1_1022<=a_1;
mulc_2_1022 : entity work.gfmul
port map(
a=>a_2,
b=>"1000000100",
X=>mulr_2_1022);

mulc_3_1022 : entity work.gfmul
port map(
a=>a_3,
b=>"0100000010",
X=>mulr_3_1022);

mulc_4_1022 : entity work.gfmul
port map(
a=>a_4,
b=>"0010000001",
X=>mulr_4_1022);

mulr_1_1023<=a_1;
mulc_2_1023 : entity work.gfmul
port map(
a=>a_2,
b=>"0000000001",
X=>mulr_2_1023);

mulc_3_1023 : entity work.gfmul
port map(
a=>a_3,
b=>"0000000001",
X=>mulr_3_1023);

mulc_4_1023 : entity work.gfmul
port map(
a=>a_4,
b=>"0000000001",
X=>mulr_4_1023);

sumr_1<= mulr_1_1 xor mulr_2_1 xor mulr_3_1 xor mulr_4_1;
sumr_2<= mulr_1_2 xor mulr_2_2 xor mulr_3_2 xor mulr_4_2;
sumr_3<= mulr_1_3 xor mulr_2_3 xor mulr_3_3 xor mulr_4_3;
sumr_4<= mulr_1_4 xor mulr_2_4 xor mulr_3_4 xor mulr_4_4;
sumr_5<= mulr_1_5 xor mulr_2_5 xor mulr_3_5 xor mulr_4_5;
sumr_6<= mulr_1_6 xor mulr_2_6 xor mulr_3_6 xor mulr_4_6;
sumr_7<= mulr_1_7 xor mulr_2_7 xor mulr_3_7 xor mulr_4_7;
sumr_8<= mulr_1_8 xor mulr_2_8 xor mulr_3_8 xor mulr_4_8;
sumr_9<= mulr_1_9 xor mulr_2_9 xor mulr_3_9 xor mulr_4_9;
sumr_10<= mulr_1_10 xor mulr_2_10 xor mulr_3_10 xor mulr_4_10;
sumr_11<= mulr_1_11 xor mulr_2_11 xor mulr_3_11 xor mulr_4_11;
sumr_12<= mulr_1_12 xor mulr_2_12 xor mulr_3_12 xor mulr_4_12;
sumr_13<= mulr_1_13 xor mulr_2_13 xor mulr_3_13 xor mulr_4_13;
sumr_14<= mulr_1_14 xor mulr_2_14 xor mulr_3_14 xor mulr_4_14;
sumr_15<= mulr_1_15 xor mulr_2_15 xor mulr_3_15 xor mulr_4_15;
sumr_16<= mulr_1_16 xor mulr_2_16 xor mulr_3_16 xor mulr_4_16;
sumr_17<= mulr_1_17 xor mulr_2_17 xor mulr_3_17 xor mulr_4_17;
sumr_18<= mulr_1_18 xor mulr_2_18 xor mulr_3_18 xor mulr_4_18;
sumr_19<= mulr_1_19 xor mulr_2_19 xor mulr_3_19 xor mulr_4_19;
sumr_20<= mulr_1_20 xor mulr_2_20 xor mulr_3_20 xor mulr_4_20;
sumr_21<= mulr_1_21 xor mulr_2_21 xor mulr_3_21 xor mulr_4_21;
sumr_22<= mulr_1_22 xor mulr_2_22 xor mulr_3_22 xor mulr_4_22;
sumr_23<= mulr_1_23 xor mulr_2_23 xor mulr_3_23 xor mulr_4_23;
sumr_24<= mulr_1_24 xor mulr_2_24 xor mulr_3_24 xor mulr_4_24;
sumr_25<= mulr_1_25 xor mulr_2_25 xor mulr_3_25 xor mulr_4_25;
sumr_26<= mulr_1_26 xor mulr_2_26 xor mulr_3_26 xor mulr_4_26;
sumr_27<= mulr_1_27 xor mulr_2_27 xor mulr_3_27 xor mulr_4_27;
sumr_28<= mulr_1_28 xor mulr_2_28 xor mulr_3_28 xor mulr_4_28;
sumr_29<= mulr_1_29 xor mulr_2_29 xor mulr_3_29 xor mulr_4_29;
sumr_30<= mulr_1_30 xor mulr_2_30 xor mulr_3_30 xor mulr_4_30;
sumr_31<= mulr_1_31 xor mulr_2_31 xor mulr_3_31 xor mulr_4_31;
sumr_32<= mulr_1_32 xor mulr_2_32 xor mulr_3_32 xor mulr_4_32;
sumr_33<= mulr_1_33 xor mulr_2_33 xor mulr_3_33 xor mulr_4_33;
sumr_34<= mulr_1_34 xor mulr_2_34 xor mulr_3_34 xor mulr_4_34;
sumr_35<= mulr_1_35 xor mulr_2_35 xor mulr_3_35 xor mulr_4_35;
sumr_36<= mulr_1_36 xor mulr_2_36 xor mulr_3_36 xor mulr_4_36;
sumr_37<= mulr_1_37 xor mulr_2_37 xor mulr_3_37 xor mulr_4_37;
sumr_38<= mulr_1_38 xor mulr_2_38 xor mulr_3_38 xor mulr_4_38;
sumr_39<= mulr_1_39 xor mulr_2_39 xor mulr_3_39 xor mulr_4_39;
sumr_40<= mulr_1_40 xor mulr_2_40 xor mulr_3_40 xor mulr_4_40;
sumr_41<= mulr_1_41 xor mulr_2_41 xor mulr_3_41 xor mulr_4_41;
sumr_42<= mulr_1_42 xor mulr_2_42 xor mulr_3_42 xor mulr_4_42;
sumr_43<= mulr_1_43 xor mulr_2_43 xor mulr_3_43 xor mulr_4_43;
sumr_44<= mulr_1_44 xor mulr_2_44 xor mulr_3_44 xor mulr_4_44;
sumr_45<= mulr_1_45 xor mulr_2_45 xor mulr_3_45 xor mulr_4_45;
sumr_46<= mulr_1_46 xor mulr_2_46 xor mulr_3_46 xor mulr_4_46;
sumr_47<= mulr_1_47 xor mulr_2_47 xor mulr_3_47 xor mulr_4_47;
sumr_48<= mulr_1_48 xor mulr_2_48 xor mulr_3_48 xor mulr_4_48;
sumr_49<= mulr_1_49 xor mulr_2_49 xor mulr_3_49 xor mulr_4_49;
sumr_50<= mulr_1_50 xor mulr_2_50 xor mulr_3_50 xor mulr_4_50;
sumr_51<= mulr_1_51 xor mulr_2_51 xor mulr_3_51 xor mulr_4_51;
sumr_52<= mulr_1_52 xor mulr_2_52 xor mulr_3_52 xor mulr_4_52;
sumr_53<= mulr_1_53 xor mulr_2_53 xor mulr_3_53 xor mulr_4_53;
sumr_54<= mulr_1_54 xor mulr_2_54 xor mulr_3_54 xor mulr_4_54;
sumr_55<= mulr_1_55 xor mulr_2_55 xor mulr_3_55 xor mulr_4_55;
sumr_56<= mulr_1_56 xor mulr_2_56 xor mulr_3_56 xor mulr_4_56;
sumr_57<= mulr_1_57 xor mulr_2_57 xor mulr_3_57 xor mulr_4_57;
sumr_58<= mulr_1_58 xor mulr_2_58 xor mulr_3_58 xor mulr_4_58;
sumr_59<= mulr_1_59 xor mulr_2_59 xor mulr_3_59 xor mulr_4_59;
sumr_60<= mulr_1_60 xor mulr_2_60 xor mulr_3_60 xor mulr_4_60;
sumr_61<= mulr_1_61 xor mulr_2_61 xor mulr_3_61 xor mulr_4_61;
sumr_62<= mulr_1_62 xor mulr_2_62 xor mulr_3_62 xor mulr_4_62;
sumr_63<= mulr_1_63 xor mulr_2_63 xor mulr_3_63 xor mulr_4_63;
sumr_64<= mulr_1_64 xor mulr_2_64 xor mulr_3_64 xor mulr_4_64;
sumr_65<= mulr_1_65 xor mulr_2_65 xor mulr_3_65 xor mulr_4_65;
sumr_66<= mulr_1_66 xor mulr_2_66 xor mulr_3_66 xor mulr_4_66;
sumr_67<= mulr_1_67 xor mulr_2_67 xor mulr_3_67 xor mulr_4_67;
sumr_68<= mulr_1_68 xor mulr_2_68 xor mulr_3_68 xor mulr_4_68;
sumr_69<= mulr_1_69 xor mulr_2_69 xor mulr_3_69 xor mulr_4_69;
sumr_70<= mulr_1_70 xor mulr_2_70 xor mulr_3_70 xor mulr_4_70;
sumr_71<= mulr_1_71 xor mulr_2_71 xor mulr_3_71 xor mulr_4_71;
sumr_72<= mulr_1_72 xor mulr_2_72 xor mulr_3_72 xor mulr_4_72;
sumr_73<= mulr_1_73 xor mulr_2_73 xor mulr_3_73 xor mulr_4_73;
sumr_74<= mulr_1_74 xor mulr_2_74 xor mulr_3_74 xor mulr_4_74;
sumr_75<= mulr_1_75 xor mulr_2_75 xor mulr_3_75 xor mulr_4_75;
sumr_76<= mulr_1_76 xor mulr_2_76 xor mulr_3_76 xor mulr_4_76;
sumr_77<= mulr_1_77 xor mulr_2_77 xor mulr_3_77 xor mulr_4_77;
sumr_78<= mulr_1_78 xor mulr_2_78 xor mulr_3_78 xor mulr_4_78;
sumr_79<= mulr_1_79 xor mulr_2_79 xor mulr_3_79 xor mulr_4_79;
sumr_80<= mulr_1_80 xor mulr_2_80 xor mulr_3_80 xor mulr_4_80;
sumr_81<= mulr_1_81 xor mulr_2_81 xor mulr_3_81 xor mulr_4_81;
sumr_82<= mulr_1_82 xor mulr_2_82 xor mulr_3_82 xor mulr_4_82;
sumr_83<= mulr_1_83 xor mulr_2_83 xor mulr_3_83 xor mulr_4_83;
sumr_84<= mulr_1_84 xor mulr_2_84 xor mulr_3_84 xor mulr_4_84;
sumr_85<= mulr_1_85 xor mulr_2_85 xor mulr_3_85 xor mulr_4_85;
sumr_86<= mulr_1_86 xor mulr_2_86 xor mulr_3_86 xor mulr_4_86;
sumr_87<= mulr_1_87 xor mulr_2_87 xor mulr_3_87 xor mulr_4_87;
sumr_88<= mulr_1_88 xor mulr_2_88 xor mulr_3_88 xor mulr_4_88;
sumr_89<= mulr_1_89 xor mulr_2_89 xor mulr_3_89 xor mulr_4_89;
sumr_90<= mulr_1_90 xor mulr_2_90 xor mulr_3_90 xor mulr_4_90;
sumr_91<= mulr_1_91 xor mulr_2_91 xor mulr_3_91 xor mulr_4_91;
sumr_92<= mulr_1_92 xor mulr_2_92 xor mulr_3_92 xor mulr_4_92;
sumr_93<= mulr_1_93 xor mulr_2_93 xor mulr_3_93 xor mulr_4_93;
sumr_94<= mulr_1_94 xor mulr_2_94 xor mulr_3_94 xor mulr_4_94;
sumr_95<= mulr_1_95 xor mulr_2_95 xor mulr_3_95 xor mulr_4_95;
sumr_96<= mulr_1_96 xor mulr_2_96 xor mulr_3_96 xor mulr_4_96;
sumr_97<= mulr_1_97 xor mulr_2_97 xor mulr_3_97 xor mulr_4_97;
sumr_98<= mulr_1_98 xor mulr_2_98 xor mulr_3_98 xor mulr_4_98;
sumr_99<= mulr_1_99 xor mulr_2_99 xor mulr_3_99 xor mulr_4_99;
sumr_100<= mulr_1_100 xor mulr_2_100 xor mulr_3_100 xor mulr_4_100;
sumr_101<= mulr_1_101 xor mulr_2_101 xor mulr_3_101 xor mulr_4_101;
sumr_102<= mulr_1_102 xor mulr_2_102 xor mulr_3_102 xor mulr_4_102;
sumr_103<= mulr_1_103 xor mulr_2_103 xor mulr_3_103 xor mulr_4_103;
sumr_104<= mulr_1_104 xor mulr_2_104 xor mulr_3_104 xor mulr_4_104;
sumr_105<= mulr_1_105 xor mulr_2_105 xor mulr_3_105 xor mulr_4_105;
sumr_106<= mulr_1_106 xor mulr_2_106 xor mulr_3_106 xor mulr_4_106;
sumr_107<= mulr_1_107 xor mulr_2_107 xor mulr_3_107 xor mulr_4_107;
sumr_108<= mulr_1_108 xor mulr_2_108 xor mulr_3_108 xor mulr_4_108;
sumr_109<= mulr_1_109 xor mulr_2_109 xor mulr_3_109 xor mulr_4_109;
sumr_110<= mulr_1_110 xor mulr_2_110 xor mulr_3_110 xor mulr_4_110;
sumr_111<= mulr_1_111 xor mulr_2_111 xor mulr_3_111 xor mulr_4_111;
sumr_112<= mulr_1_112 xor mulr_2_112 xor mulr_3_112 xor mulr_4_112;
sumr_113<= mulr_1_113 xor mulr_2_113 xor mulr_3_113 xor mulr_4_113;
sumr_114<= mulr_1_114 xor mulr_2_114 xor mulr_3_114 xor mulr_4_114;
sumr_115<= mulr_1_115 xor mulr_2_115 xor mulr_3_115 xor mulr_4_115;
sumr_116<= mulr_1_116 xor mulr_2_116 xor mulr_3_116 xor mulr_4_116;
sumr_117<= mulr_1_117 xor mulr_2_117 xor mulr_3_117 xor mulr_4_117;
sumr_118<= mulr_1_118 xor mulr_2_118 xor mulr_3_118 xor mulr_4_118;
sumr_119<= mulr_1_119 xor mulr_2_119 xor mulr_3_119 xor mulr_4_119;
sumr_120<= mulr_1_120 xor mulr_2_120 xor mulr_3_120 xor mulr_4_120;
sumr_121<= mulr_1_121 xor mulr_2_121 xor mulr_3_121 xor mulr_4_121;
sumr_122<= mulr_1_122 xor mulr_2_122 xor mulr_3_122 xor mulr_4_122;
sumr_123<= mulr_1_123 xor mulr_2_123 xor mulr_3_123 xor mulr_4_123;
sumr_124<= mulr_1_124 xor mulr_2_124 xor mulr_3_124 xor mulr_4_124;
sumr_125<= mulr_1_125 xor mulr_2_125 xor mulr_3_125 xor mulr_4_125;
sumr_126<= mulr_1_126 xor mulr_2_126 xor mulr_3_126 xor mulr_4_126;
sumr_127<= mulr_1_127 xor mulr_2_127 xor mulr_3_127 xor mulr_4_127;
sumr_128<= mulr_1_128 xor mulr_2_128 xor mulr_3_128 xor mulr_4_128;
sumr_129<= mulr_1_129 xor mulr_2_129 xor mulr_3_129 xor mulr_4_129;
sumr_130<= mulr_1_130 xor mulr_2_130 xor mulr_3_130 xor mulr_4_130;
sumr_131<= mulr_1_131 xor mulr_2_131 xor mulr_3_131 xor mulr_4_131;
sumr_132<= mulr_1_132 xor mulr_2_132 xor mulr_3_132 xor mulr_4_132;
sumr_133<= mulr_1_133 xor mulr_2_133 xor mulr_3_133 xor mulr_4_133;
sumr_134<= mulr_1_134 xor mulr_2_134 xor mulr_3_134 xor mulr_4_134;
sumr_135<= mulr_1_135 xor mulr_2_135 xor mulr_3_135 xor mulr_4_135;
sumr_136<= mulr_1_136 xor mulr_2_136 xor mulr_3_136 xor mulr_4_136;
sumr_137<= mulr_1_137 xor mulr_2_137 xor mulr_3_137 xor mulr_4_137;
sumr_138<= mulr_1_138 xor mulr_2_138 xor mulr_3_138 xor mulr_4_138;
sumr_139<= mulr_1_139 xor mulr_2_139 xor mulr_3_139 xor mulr_4_139;
sumr_140<= mulr_1_140 xor mulr_2_140 xor mulr_3_140 xor mulr_4_140;
sumr_141<= mulr_1_141 xor mulr_2_141 xor mulr_3_141 xor mulr_4_141;
sumr_142<= mulr_1_142 xor mulr_2_142 xor mulr_3_142 xor mulr_4_142;
sumr_143<= mulr_1_143 xor mulr_2_143 xor mulr_3_143 xor mulr_4_143;
sumr_144<= mulr_1_144 xor mulr_2_144 xor mulr_3_144 xor mulr_4_144;
sumr_145<= mulr_1_145 xor mulr_2_145 xor mulr_3_145 xor mulr_4_145;
sumr_146<= mulr_1_146 xor mulr_2_146 xor mulr_3_146 xor mulr_4_146;
sumr_147<= mulr_1_147 xor mulr_2_147 xor mulr_3_147 xor mulr_4_147;
sumr_148<= mulr_1_148 xor mulr_2_148 xor mulr_3_148 xor mulr_4_148;
sumr_149<= mulr_1_149 xor mulr_2_149 xor mulr_3_149 xor mulr_4_149;
sumr_150<= mulr_1_150 xor mulr_2_150 xor mulr_3_150 xor mulr_4_150;
sumr_151<= mulr_1_151 xor mulr_2_151 xor mulr_3_151 xor mulr_4_151;
sumr_152<= mulr_1_152 xor mulr_2_152 xor mulr_3_152 xor mulr_4_152;
sumr_153<= mulr_1_153 xor mulr_2_153 xor mulr_3_153 xor mulr_4_153;
sumr_154<= mulr_1_154 xor mulr_2_154 xor mulr_3_154 xor mulr_4_154;
sumr_155<= mulr_1_155 xor mulr_2_155 xor mulr_3_155 xor mulr_4_155;
sumr_156<= mulr_1_156 xor mulr_2_156 xor mulr_3_156 xor mulr_4_156;
sumr_157<= mulr_1_157 xor mulr_2_157 xor mulr_3_157 xor mulr_4_157;
sumr_158<= mulr_1_158 xor mulr_2_158 xor mulr_3_158 xor mulr_4_158;
sumr_159<= mulr_1_159 xor mulr_2_159 xor mulr_3_159 xor mulr_4_159;
sumr_160<= mulr_1_160 xor mulr_2_160 xor mulr_3_160 xor mulr_4_160;
sumr_161<= mulr_1_161 xor mulr_2_161 xor mulr_3_161 xor mulr_4_161;
sumr_162<= mulr_1_162 xor mulr_2_162 xor mulr_3_162 xor mulr_4_162;
sumr_163<= mulr_1_163 xor mulr_2_163 xor mulr_3_163 xor mulr_4_163;
sumr_164<= mulr_1_164 xor mulr_2_164 xor mulr_3_164 xor mulr_4_164;
sumr_165<= mulr_1_165 xor mulr_2_165 xor mulr_3_165 xor mulr_4_165;
sumr_166<= mulr_1_166 xor mulr_2_166 xor mulr_3_166 xor mulr_4_166;
sumr_167<= mulr_1_167 xor mulr_2_167 xor mulr_3_167 xor mulr_4_167;
sumr_168<= mulr_1_168 xor mulr_2_168 xor mulr_3_168 xor mulr_4_168;
sumr_169<= mulr_1_169 xor mulr_2_169 xor mulr_3_169 xor mulr_4_169;
sumr_170<= mulr_1_170 xor mulr_2_170 xor mulr_3_170 xor mulr_4_170;
sumr_171<= mulr_1_171 xor mulr_2_171 xor mulr_3_171 xor mulr_4_171;
sumr_172<= mulr_1_172 xor mulr_2_172 xor mulr_3_172 xor mulr_4_172;
sumr_173<= mulr_1_173 xor mulr_2_173 xor mulr_3_173 xor mulr_4_173;
sumr_174<= mulr_1_174 xor mulr_2_174 xor mulr_3_174 xor mulr_4_174;
sumr_175<= mulr_1_175 xor mulr_2_175 xor mulr_3_175 xor mulr_4_175;
sumr_176<= mulr_1_176 xor mulr_2_176 xor mulr_3_176 xor mulr_4_176;
sumr_177<= mulr_1_177 xor mulr_2_177 xor mulr_3_177 xor mulr_4_177;
sumr_178<= mulr_1_178 xor mulr_2_178 xor mulr_3_178 xor mulr_4_178;
sumr_179<= mulr_1_179 xor mulr_2_179 xor mulr_3_179 xor mulr_4_179;
sumr_180<= mulr_1_180 xor mulr_2_180 xor mulr_3_180 xor mulr_4_180;
sumr_181<= mulr_1_181 xor mulr_2_181 xor mulr_3_181 xor mulr_4_181;
sumr_182<= mulr_1_182 xor mulr_2_182 xor mulr_3_182 xor mulr_4_182;
sumr_183<= mulr_1_183 xor mulr_2_183 xor mulr_3_183 xor mulr_4_183;
sumr_184<= mulr_1_184 xor mulr_2_184 xor mulr_3_184 xor mulr_4_184;
sumr_185<= mulr_1_185 xor mulr_2_185 xor mulr_3_185 xor mulr_4_185;
sumr_186<= mulr_1_186 xor mulr_2_186 xor mulr_3_186 xor mulr_4_186;
sumr_187<= mulr_1_187 xor mulr_2_187 xor mulr_3_187 xor mulr_4_187;
sumr_188<= mulr_1_188 xor mulr_2_188 xor mulr_3_188 xor mulr_4_188;
sumr_189<= mulr_1_189 xor mulr_2_189 xor mulr_3_189 xor mulr_4_189;
sumr_190<= mulr_1_190 xor mulr_2_190 xor mulr_3_190 xor mulr_4_190;
sumr_191<= mulr_1_191 xor mulr_2_191 xor mulr_3_191 xor mulr_4_191;
sumr_192<= mulr_1_192 xor mulr_2_192 xor mulr_3_192 xor mulr_4_192;
sumr_193<= mulr_1_193 xor mulr_2_193 xor mulr_3_193 xor mulr_4_193;
sumr_194<= mulr_1_194 xor mulr_2_194 xor mulr_3_194 xor mulr_4_194;
sumr_195<= mulr_1_195 xor mulr_2_195 xor mulr_3_195 xor mulr_4_195;
sumr_196<= mulr_1_196 xor mulr_2_196 xor mulr_3_196 xor mulr_4_196;
sumr_197<= mulr_1_197 xor mulr_2_197 xor mulr_3_197 xor mulr_4_197;
sumr_198<= mulr_1_198 xor mulr_2_198 xor mulr_3_198 xor mulr_4_198;
sumr_199<= mulr_1_199 xor mulr_2_199 xor mulr_3_199 xor mulr_4_199;
sumr_200<= mulr_1_200 xor mulr_2_200 xor mulr_3_200 xor mulr_4_200;
sumr_201<= mulr_1_201 xor mulr_2_201 xor mulr_3_201 xor mulr_4_201;
sumr_202<= mulr_1_202 xor mulr_2_202 xor mulr_3_202 xor mulr_4_202;
sumr_203<= mulr_1_203 xor mulr_2_203 xor mulr_3_203 xor mulr_4_203;
sumr_204<= mulr_1_204 xor mulr_2_204 xor mulr_3_204 xor mulr_4_204;
sumr_205<= mulr_1_205 xor mulr_2_205 xor mulr_3_205 xor mulr_4_205;
sumr_206<= mulr_1_206 xor mulr_2_206 xor mulr_3_206 xor mulr_4_206;
sumr_207<= mulr_1_207 xor mulr_2_207 xor mulr_3_207 xor mulr_4_207;
sumr_208<= mulr_1_208 xor mulr_2_208 xor mulr_3_208 xor mulr_4_208;
sumr_209<= mulr_1_209 xor mulr_2_209 xor mulr_3_209 xor mulr_4_209;
sumr_210<= mulr_1_210 xor mulr_2_210 xor mulr_3_210 xor mulr_4_210;
sumr_211<= mulr_1_211 xor mulr_2_211 xor mulr_3_211 xor mulr_4_211;
sumr_212<= mulr_1_212 xor mulr_2_212 xor mulr_3_212 xor mulr_4_212;
sumr_213<= mulr_1_213 xor mulr_2_213 xor mulr_3_213 xor mulr_4_213;
sumr_214<= mulr_1_214 xor mulr_2_214 xor mulr_3_214 xor mulr_4_214;
sumr_215<= mulr_1_215 xor mulr_2_215 xor mulr_3_215 xor mulr_4_215;
sumr_216<= mulr_1_216 xor mulr_2_216 xor mulr_3_216 xor mulr_4_216;
sumr_217<= mulr_1_217 xor mulr_2_217 xor mulr_3_217 xor mulr_4_217;
sumr_218<= mulr_1_218 xor mulr_2_218 xor mulr_3_218 xor mulr_4_218;
sumr_219<= mulr_1_219 xor mulr_2_219 xor mulr_3_219 xor mulr_4_219;
sumr_220<= mulr_1_220 xor mulr_2_220 xor mulr_3_220 xor mulr_4_220;
sumr_221<= mulr_1_221 xor mulr_2_221 xor mulr_3_221 xor mulr_4_221;
sumr_222<= mulr_1_222 xor mulr_2_222 xor mulr_3_222 xor mulr_4_222;
sumr_223<= mulr_1_223 xor mulr_2_223 xor mulr_3_223 xor mulr_4_223;
sumr_224<= mulr_1_224 xor mulr_2_224 xor mulr_3_224 xor mulr_4_224;
sumr_225<= mulr_1_225 xor mulr_2_225 xor mulr_3_225 xor mulr_4_225;
sumr_226<= mulr_1_226 xor mulr_2_226 xor mulr_3_226 xor mulr_4_226;
sumr_227<= mulr_1_227 xor mulr_2_227 xor mulr_3_227 xor mulr_4_227;
sumr_228<= mulr_1_228 xor mulr_2_228 xor mulr_3_228 xor mulr_4_228;
sumr_229<= mulr_1_229 xor mulr_2_229 xor mulr_3_229 xor mulr_4_229;
sumr_230<= mulr_1_230 xor mulr_2_230 xor mulr_3_230 xor mulr_4_230;
sumr_231<= mulr_1_231 xor mulr_2_231 xor mulr_3_231 xor mulr_4_231;
sumr_232<= mulr_1_232 xor mulr_2_232 xor mulr_3_232 xor mulr_4_232;
sumr_233<= mulr_1_233 xor mulr_2_233 xor mulr_3_233 xor mulr_4_233;
sumr_234<= mulr_1_234 xor mulr_2_234 xor mulr_3_234 xor mulr_4_234;
sumr_235<= mulr_1_235 xor mulr_2_235 xor mulr_3_235 xor mulr_4_235;
sumr_236<= mulr_1_236 xor mulr_2_236 xor mulr_3_236 xor mulr_4_236;
sumr_237<= mulr_1_237 xor mulr_2_237 xor mulr_3_237 xor mulr_4_237;
sumr_238<= mulr_1_238 xor mulr_2_238 xor mulr_3_238 xor mulr_4_238;
sumr_239<= mulr_1_239 xor mulr_2_239 xor mulr_3_239 xor mulr_4_239;
sumr_240<= mulr_1_240 xor mulr_2_240 xor mulr_3_240 xor mulr_4_240;
sumr_241<= mulr_1_241 xor mulr_2_241 xor mulr_3_241 xor mulr_4_241;
sumr_242<= mulr_1_242 xor mulr_2_242 xor mulr_3_242 xor mulr_4_242;
sumr_243<= mulr_1_243 xor mulr_2_243 xor mulr_3_243 xor mulr_4_243;
sumr_244<= mulr_1_244 xor mulr_2_244 xor mulr_3_244 xor mulr_4_244;
sumr_245<= mulr_1_245 xor mulr_2_245 xor mulr_3_245 xor mulr_4_245;
sumr_246<= mulr_1_246 xor mulr_2_246 xor mulr_3_246 xor mulr_4_246;
sumr_247<= mulr_1_247 xor mulr_2_247 xor mulr_3_247 xor mulr_4_247;
sumr_248<= mulr_1_248 xor mulr_2_248 xor mulr_3_248 xor mulr_4_248;
sumr_249<= mulr_1_249 xor mulr_2_249 xor mulr_3_249 xor mulr_4_249;
sumr_250<= mulr_1_250 xor mulr_2_250 xor mulr_3_250 xor mulr_4_250;
sumr_251<= mulr_1_251 xor mulr_2_251 xor mulr_3_251 xor mulr_4_251;
sumr_252<= mulr_1_252 xor mulr_2_252 xor mulr_3_252 xor mulr_4_252;
sumr_253<= mulr_1_253 xor mulr_2_253 xor mulr_3_253 xor mulr_4_253;
sumr_254<= mulr_1_254 xor mulr_2_254 xor mulr_3_254 xor mulr_4_254;
sumr_255<= mulr_1_255 xor mulr_2_255 xor mulr_3_255 xor mulr_4_255;
sumr_256<= mulr_1_256 xor mulr_2_256 xor mulr_3_256 xor mulr_4_256;
sumr_257<= mulr_1_257 xor mulr_2_257 xor mulr_3_257 xor mulr_4_257;
sumr_258<= mulr_1_258 xor mulr_2_258 xor mulr_3_258 xor mulr_4_258;
sumr_259<= mulr_1_259 xor mulr_2_259 xor mulr_3_259 xor mulr_4_259;
sumr_260<= mulr_1_260 xor mulr_2_260 xor mulr_3_260 xor mulr_4_260;
sumr_261<= mulr_1_261 xor mulr_2_261 xor mulr_3_261 xor mulr_4_261;
sumr_262<= mulr_1_262 xor mulr_2_262 xor mulr_3_262 xor mulr_4_262;
sumr_263<= mulr_1_263 xor mulr_2_263 xor mulr_3_263 xor mulr_4_263;
sumr_264<= mulr_1_264 xor mulr_2_264 xor mulr_3_264 xor mulr_4_264;
sumr_265<= mulr_1_265 xor mulr_2_265 xor mulr_3_265 xor mulr_4_265;
sumr_266<= mulr_1_266 xor mulr_2_266 xor mulr_3_266 xor mulr_4_266;
sumr_267<= mulr_1_267 xor mulr_2_267 xor mulr_3_267 xor mulr_4_267;
sumr_268<= mulr_1_268 xor mulr_2_268 xor mulr_3_268 xor mulr_4_268;
sumr_269<= mulr_1_269 xor mulr_2_269 xor mulr_3_269 xor mulr_4_269;
sumr_270<= mulr_1_270 xor mulr_2_270 xor mulr_3_270 xor mulr_4_270;
sumr_271<= mulr_1_271 xor mulr_2_271 xor mulr_3_271 xor mulr_4_271;
sumr_272<= mulr_1_272 xor mulr_2_272 xor mulr_3_272 xor mulr_4_272;
sumr_273<= mulr_1_273 xor mulr_2_273 xor mulr_3_273 xor mulr_4_273;
sumr_274<= mulr_1_274 xor mulr_2_274 xor mulr_3_274 xor mulr_4_274;
sumr_275<= mulr_1_275 xor mulr_2_275 xor mulr_3_275 xor mulr_4_275;
sumr_276<= mulr_1_276 xor mulr_2_276 xor mulr_3_276 xor mulr_4_276;
sumr_277<= mulr_1_277 xor mulr_2_277 xor mulr_3_277 xor mulr_4_277;
sumr_278<= mulr_1_278 xor mulr_2_278 xor mulr_3_278 xor mulr_4_278;
sumr_279<= mulr_1_279 xor mulr_2_279 xor mulr_3_279 xor mulr_4_279;
sumr_280<= mulr_1_280 xor mulr_2_280 xor mulr_3_280 xor mulr_4_280;
sumr_281<= mulr_1_281 xor mulr_2_281 xor mulr_3_281 xor mulr_4_281;
sumr_282<= mulr_1_282 xor mulr_2_282 xor mulr_3_282 xor mulr_4_282;
sumr_283<= mulr_1_283 xor mulr_2_283 xor mulr_3_283 xor mulr_4_283;
sumr_284<= mulr_1_284 xor mulr_2_284 xor mulr_3_284 xor mulr_4_284;
sumr_285<= mulr_1_285 xor mulr_2_285 xor mulr_3_285 xor mulr_4_285;
sumr_286<= mulr_1_286 xor mulr_2_286 xor mulr_3_286 xor mulr_4_286;
sumr_287<= mulr_1_287 xor mulr_2_287 xor mulr_3_287 xor mulr_4_287;
sumr_288<= mulr_1_288 xor mulr_2_288 xor mulr_3_288 xor mulr_4_288;
sumr_289<= mulr_1_289 xor mulr_2_289 xor mulr_3_289 xor mulr_4_289;
sumr_290<= mulr_1_290 xor mulr_2_290 xor mulr_3_290 xor mulr_4_290;
sumr_291<= mulr_1_291 xor mulr_2_291 xor mulr_3_291 xor mulr_4_291;
sumr_292<= mulr_1_292 xor mulr_2_292 xor mulr_3_292 xor mulr_4_292;
sumr_293<= mulr_1_293 xor mulr_2_293 xor mulr_3_293 xor mulr_4_293;
sumr_294<= mulr_1_294 xor mulr_2_294 xor mulr_3_294 xor mulr_4_294;
sumr_295<= mulr_1_295 xor mulr_2_295 xor mulr_3_295 xor mulr_4_295;
sumr_296<= mulr_1_296 xor mulr_2_296 xor mulr_3_296 xor mulr_4_296;
sumr_297<= mulr_1_297 xor mulr_2_297 xor mulr_3_297 xor mulr_4_297;
sumr_298<= mulr_1_298 xor mulr_2_298 xor mulr_3_298 xor mulr_4_298;
sumr_299<= mulr_1_299 xor mulr_2_299 xor mulr_3_299 xor mulr_4_299;
sumr_300<= mulr_1_300 xor mulr_2_300 xor mulr_3_300 xor mulr_4_300;
sumr_301<= mulr_1_301 xor mulr_2_301 xor mulr_3_301 xor mulr_4_301;
sumr_302<= mulr_1_302 xor mulr_2_302 xor mulr_3_302 xor mulr_4_302;
sumr_303<= mulr_1_303 xor mulr_2_303 xor mulr_3_303 xor mulr_4_303;
sumr_304<= mulr_1_304 xor mulr_2_304 xor mulr_3_304 xor mulr_4_304;
sumr_305<= mulr_1_305 xor mulr_2_305 xor mulr_3_305 xor mulr_4_305;
sumr_306<= mulr_1_306 xor mulr_2_306 xor mulr_3_306 xor mulr_4_306;
sumr_307<= mulr_1_307 xor mulr_2_307 xor mulr_3_307 xor mulr_4_307;
sumr_308<= mulr_1_308 xor mulr_2_308 xor mulr_3_308 xor mulr_4_308;
sumr_309<= mulr_1_309 xor mulr_2_309 xor mulr_3_309 xor mulr_4_309;
sumr_310<= mulr_1_310 xor mulr_2_310 xor mulr_3_310 xor mulr_4_310;
sumr_311<= mulr_1_311 xor mulr_2_311 xor mulr_3_311 xor mulr_4_311;
sumr_312<= mulr_1_312 xor mulr_2_312 xor mulr_3_312 xor mulr_4_312;
sumr_313<= mulr_1_313 xor mulr_2_313 xor mulr_3_313 xor mulr_4_313;
sumr_314<= mulr_1_314 xor mulr_2_314 xor mulr_3_314 xor mulr_4_314;
sumr_315<= mulr_1_315 xor mulr_2_315 xor mulr_3_315 xor mulr_4_315;
sumr_316<= mulr_1_316 xor mulr_2_316 xor mulr_3_316 xor mulr_4_316;
sumr_317<= mulr_1_317 xor mulr_2_317 xor mulr_3_317 xor mulr_4_317;
sumr_318<= mulr_1_318 xor mulr_2_318 xor mulr_3_318 xor mulr_4_318;
sumr_319<= mulr_1_319 xor mulr_2_319 xor mulr_3_319 xor mulr_4_319;
sumr_320<= mulr_1_320 xor mulr_2_320 xor mulr_3_320 xor mulr_4_320;
sumr_321<= mulr_1_321 xor mulr_2_321 xor mulr_3_321 xor mulr_4_321;
sumr_322<= mulr_1_322 xor mulr_2_322 xor mulr_3_322 xor mulr_4_322;
sumr_323<= mulr_1_323 xor mulr_2_323 xor mulr_3_323 xor mulr_4_323;
sumr_324<= mulr_1_324 xor mulr_2_324 xor mulr_3_324 xor mulr_4_324;
sumr_325<= mulr_1_325 xor mulr_2_325 xor mulr_3_325 xor mulr_4_325;
sumr_326<= mulr_1_326 xor mulr_2_326 xor mulr_3_326 xor mulr_4_326;
sumr_327<= mulr_1_327 xor mulr_2_327 xor mulr_3_327 xor mulr_4_327;
sumr_328<= mulr_1_328 xor mulr_2_328 xor mulr_3_328 xor mulr_4_328;
sumr_329<= mulr_1_329 xor mulr_2_329 xor mulr_3_329 xor mulr_4_329;
sumr_330<= mulr_1_330 xor mulr_2_330 xor mulr_3_330 xor mulr_4_330;
sumr_331<= mulr_1_331 xor mulr_2_331 xor mulr_3_331 xor mulr_4_331;
sumr_332<= mulr_1_332 xor mulr_2_332 xor mulr_3_332 xor mulr_4_332;
sumr_333<= mulr_1_333 xor mulr_2_333 xor mulr_3_333 xor mulr_4_333;
sumr_334<= mulr_1_334 xor mulr_2_334 xor mulr_3_334 xor mulr_4_334;
sumr_335<= mulr_1_335 xor mulr_2_335 xor mulr_3_335 xor mulr_4_335;
sumr_336<= mulr_1_336 xor mulr_2_336 xor mulr_3_336 xor mulr_4_336;
sumr_337<= mulr_1_337 xor mulr_2_337 xor mulr_3_337 xor mulr_4_337;
sumr_338<= mulr_1_338 xor mulr_2_338 xor mulr_3_338 xor mulr_4_338;
sumr_339<= mulr_1_339 xor mulr_2_339 xor mulr_3_339 xor mulr_4_339;
sumr_340<= mulr_1_340 xor mulr_2_340 xor mulr_3_340 xor mulr_4_340;
sumr_341<= mulr_1_341 xor mulr_2_341 xor mulr_3_341 xor mulr_4_341;
sumr_342<= mulr_1_342 xor mulr_2_342 xor mulr_3_342 xor mulr_4_342;
sumr_343<= mulr_1_343 xor mulr_2_343 xor mulr_3_343 xor mulr_4_343;
sumr_344<= mulr_1_344 xor mulr_2_344 xor mulr_3_344 xor mulr_4_344;
sumr_345<= mulr_1_345 xor mulr_2_345 xor mulr_3_345 xor mulr_4_345;
sumr_346<= mulr_1_346 xor mulr_2_346 xor mulr_3_346 xor mulr_4_346;
sumr_347<= mulr_1_347 xor mulr_2_347 xor mulr_3_347 xor mulr_4_347;
sumr_348<= mulr_1_348 xor mulr_2_348 xor mulr_3_348 xor mulr_4_348;
sumr_349<= mulr_1_349 xor mulr_2_349 xor mulr_3_349 xor mulr_4_349;
sumr_350<= mulr_1_350 xor mulr_2_350 xor mulr_3_350 xor mulr_4_350;
sumr_351<= mulr_1_351 xor mulr_2_351 xor mulr_3_351 xor mulr_4_351;
sumr_352<= mulr_1_352 xor mulr_2_352 xor mulr_3_352 xor mulr_4_352;
sumr_353<= mulr_1_353 xor mulr_2_353 xor mulr_3_353 xor mulr_4_353;
sumr_354<= mulr_1_354 xor mulr_2_354 xor mulr_3_354 xor mulr_4_354;
sumr_355<= mulr_1_355 xor mulr_2_355 xor mulr_3_355 xor mulr_4_355;
sumr_356<= mulr_1_356 xor mulr_2_356 xor mulr_3_356 xor mulr_4_356;
sumr_357<= mulr_1_357 xor mulr_2_357 xor mulr_3_357 xor mulr_4_357;
sumr_358<= mulr_1_358 xor mulr_2_358 xor mulr_3_358 xor mulr_4_358;
sumr_359<= mulr_1_359 xor mulr_2_359 xor mulr_3_359 xor mulr_4_359;
sumr_360<= mulr_1_360 xor mulr_2_360 xor mulr_3_360 xor mulr_4_360;
sumr_361<= mulr_1_361 xor mulr_2_361 xor mulr_3_361 xor mulr_4_361;
sumr_362<= mulr_1_362 xor mulr_2_362 xor mulr_3_362 xor mulr_4_362;
sumr_363<= mulr_1_363 xor mulr_2_363 xor mulr_3_363 xor mulr_4_363;
sumr_364<= mulr_1_364 xor mulr_2_364 xor mulr_3_364 xor mulr_4_364;
sumr_365<= mulr_1_365 xor mulr_2_365 xor mulr_3_365 xor mulr_4_365;
sumr_366<= mulr_1_366 xor mulr_2_366 xor mulr_3_366 xor mulr_4_366;
sumr_367<= mulr_1_367 xor mulr_2_367 xor mulr_3_367 xor mulr_4_367;
sumr_368<= mulr_1_368 xor mulr_2_368 xor mulr_3_368 xor mulr_4_368;
sumr_369<= mulr_1_369 xor mulr_2_369 xor mulr_3_369 xor mulr_4_369;
sumr_370<= mulr_1_370 xor mulr_2_370 xor mulr_3_370 xor mulr_4_370;
sumr_371<= mulr_1_371 xor mulr_2_371 xor mulr_3_371 xor mulr_4_371;
sumr_372<= mulr_1_372 xor mulr_2_372 xor mulr_3_372 xor mulr_4_372;
sumr_373<= mulr_1_373 xor mulr_2_373 xor mulr_3_373 xor mulr_4_373;
sumr_374<= mulr_1_374 xor mulr_2_374 xor mulr_3_374 xor mulr_4_374;
sumr_375<= mulr_1_375 xor mulr_2_375 xor mulr_3_375 xor mulr_4_375;
sumr_376<= mulr_1_376 xor mulr_2_376 xor mulr_3_376 xor mulr_4_376;
sumr_377<= mulr_1_377 xor mulr_2_377 xor mulr_3_377 xor mulr_4_377;
sumr_378<= mulr_1_378 xor mulr_2_378 xor mulr_3_378 xor mulr_4_378;
sumr_379<= mulr_1_379 xor mulr_2_379 xor mulr_3_379 xor mulr_4_379;
sumr_380<= mulr_1_380 xor mulr_2_380 xor mulr_3_380 xor mulr_4_380;
sumr_381<= mulr_1_381 xor mulr_2_381 xor mulr_3_381 xor mulr_4_381;
sumr_382<= mulr_1_382 xor mulr_2_382 xor mulr_3_382 xor mulr_4_382;
sumr_383<= mulr_1_383 xor mulr_2_383 xor mulr_3_383 xor mulr_4_383;
sumr_384<= mulr_1_384 xor mulr_2_384 xor mulr_3_384 xor mulr_4_384;
sumr_385<= mulr_1_385 xor mulr_2_385 xor mulr_3_385 xor mulr_4_385;
sumr_386<= mulr_1_386 xor mulr_2_386 xor mulr_3_386 xor mulr_4_386;
sumr_387<= mulr_1_387 xor mulr_2_387 xor mulr_3_387 xor mulr_4_387;
sumr_388<= mulr_1_388 xor mulr_2_388 xor mulr_3_388 xor mulr_4_388;
sumr_389<= mulr_1_389 xor mulr_2_389 xor mulr_3_389 xor mulr_4_389;
sumr_390<= mulr_1_390 xor mulr_2_390 xor mulr_3_390 xor mulr_4_390;
sumr_391<= mulr_1_391 xor mulr_2_391 xor mulr_3_391 xor mulr_4_391;
sumr_392<= mulr_1_392 xor mulr_2_392 xor mulr_3_392 xor mulr_4_392;
sumr_393<= mulr_1_393 xor mulr_2_393 xor mulr_3_393 xor mulr_4_393;
sumr_394<= mulr_1_394 xor mulr_2_394 xor mulr_3_394 xor mulr_4_394;
sumr_395<= mulr_1_395 xor mulr_2_395 xor mulr_3_395 xor mulr_4_395;
sumr_396<= mulr_1_396 xor mulr_2_396 xor mulr_3_396 xor mulr_4_396;
sumr_397<= mulr_1_397 xor mulr_2_397 xor mulr_3_397 xor mulr_4_397;
sumr_398<= mulr_1_398 xor mulr_2_398 xor mulr_3_398 xor mulr_4_398;
sumr_399<= mulr_1_399 xor mulr_2_399 xor mulr_3_399 xor mulr_4_399;
sumr_400<= mulr_1_400 xor mulr_2_400 xor mulr_3_400 xor mulr_4_400;
sumr_401<= mulr_1_401 xor mulr_2_401 xor mulr_3_401 xor mulr_4_401;
sumr_402<= mulr_1_402 xor mulr_2_402 xor mulr_3_402 xor mulr_4_402;
sumr_403<= mulr_1_403 xor mulr_2_403 xor mulr_3_403 xor mulr_4_403;
sumr_404<= mulr_1_404 xor mulr_2_404 xor mulr_3_404 xor mulr_4_404;
sumr_405<= mulr_1_405 xor mulr_2_405 xor mulr_3_405 xor mulr_4_405;
sumr_406<= mulr_1_406 xor mulr_2_406 xor mulr_3_406 xor mulr_4_406;
sumr_407<= mulr_1_407 xor mulr_2_407 xor mulr_3_407 xor mulr_4_407;
sumr_408<= mulr_1_408 xor mulr_2_408 xor mulr_3_408 xor mulr_4_408;
sumr_409<= mulr_1_409 xor mulr_2_409 xor mulr_3_409 xor mulr_4_409;
sumr_410<= mulr_1_410 xor mulr_2_410 xor mulr_3_410 xor mulr_4_410;
sumr_411<= mulr_1_411 xor mulr_2_411 xor mulr_3_411 xor mulr_4_411;
sumr_412<= mulr_1_412 xor mulr_2_412 xor mulr_3_412 xor mulr_4_412;
sumr_413<= mulr_1_413 xor mulr_2_413 xor mulr_3_413 xor mulr_4_413;
sumr_414<= mulr_1_414 xor mulr_2_414 xor mulr_3_414 xor mulr_4_414;
sumr_415<= mulr_1_415 xor mulr_2_415 xor mulr_3_415 xor mulr_4_415;
sumr_416<= mulr_1_416 xor mulr_2_416 xor mulr_3_416 xor mulr_4_416;
sumr_417<= mulr_1_417 xor mulr_2_417 xor mulr_3_417 xor mulr_4_417;
sumr_418<= mulr_1_418 xor mulr_2_418 xor mulr_3_418 xor mulr_4_418;
sumr_419<= mulr_1_419 xor mulr_2_419 xor mulr_3_419 xor mulr_4_419;
sumr_420<= mulr_1_420 xor mulr_2_420 xor mulr_3_420 xor mulr_4_420;
sumr_421<= mulr_1_421 xor mulr_2_421 xor mulr_3_421 xor mulr_4_421;
sumr_422<= mulr_1_422 xor mulr_2_422 xor mulr_3_422 xor mulr_4_422;
sumr_423<= mulr_1_423 xor mulr_2_423 xor mulr_3_423 xor mulr_4_423;
sumr_424<= mulr_1_424 xor mulr_2_424 xor mulr_3_424 xor mulr_4_424;
sumr_425<= mulr_1_425 xor mulr_2_425 xor mulr_3_425 xor mulr_4_425;
sumr_426<= mulr_1_426 xor mulr_2_426 xor mulr_3_426 xor mulr_4_426;
sumr_427<= mulr_1_427 xor mulr_2_427 xor mulr_3_427 xor mulr_4_427;
sumr_428<= mulr_1_428 xor mulr_2_428 xor mulr_3_428 xor mulr_4_428;
sumr_429<= mulr_1_429 xor mulr_2_429 xor mulr_3_429 xor mulr_4_429;
sumr_430<= mulr_1_430 xor mulr_2_430 xor mulr_3_430 xor mulr_4_430;
sumr_431<= mulr_1_431 xor mulr_2_431 xor mulr_3_431 xor mulr_4_431;
sumr_432<= mulr_1_432 xor mulr_2_432 xor mulr_3_432 xor mulr_4_432;
sumr_433<= mulr_1_433 xor mulr_2_433 xor mulr_3_433 xor mulr_4_433;
sumr_434<= mulr_1_434 xor mulr_2_434 xor mulr_3_434 xor mulr_4_434;
sumr_435<= mulr_1_435 xor mulr_2_435 xor mulr_3_435 xor mulr_4_435;
sumr_436<= mulr_1_436 xor mulr_2_436 xor mulr_3_436 xor mulr_4_436;
sumr_437<= mulr_1_437 xor mulr_2_437 xor mulr_3_437 xor mulr_4_437;
sumr_438<= mulr_1_438 xor mulr_2_438 xor mulr_3_438 xor mulr_4_438;
sumr_439<= mulr_1_439 xor mulr_2_439 xor mulr_3_439 xor mulr_4_439;
sumr_440<= mulr_1_440 xor mulr_2_440 xor mulr_3_440 xor mulr_4_440;
sumr_441<= mulr_1_441 xor mulr_2_441 xor mulr_3_441 xor mulr_4_441;
sumr_442<= mulr_1_442 xor mulr_2_442 xor mulr_3_442 xor mulr_4_442;
sumr_443<= mulr_1_443 xor mulr_2_443 xor mulr_3_443 xor mulr_4_443;
sumr_444<= mulr_1_444 xor mulr_2_444 xor mulr_3_444 xor mulr_4_444;
sumr_445<= mulr_1_445 xor mulr_2_445 xor mulr_3_445 xor mulr_4_445;
sumr_446<= mulr_1_446 xor mulr_2_446 xor mulr_3_446 xor mulr_4_446;
sumr_447<= mulr_1_447 xor mulr_2_447 xor mulr_3_447 xor mulr_4_447;
sumr_448<= mulr_1_448 xor mulr_2_448 xor mulr_3_448 xor mulr_4_448;
sumr_449<= mulr_1_449 xor mulr_2_449 xor mulr_3_449 xor mulr_4_449;
sumr_450<= mulr_1_450 xor mulr_2_450 xor mulr_3_450 xor mulr_4_450;
sumr_451<= mulr_1_451 xor mulr_2_451 xor mulr_3_451 xor mulr_4_451;
sumr_452<= mulr_1_452 xor mulr_2_452 xor mulr_3_452 xor mulr_4_452;
sumr_453<= mulr_1_453 xor mulr_2_453 xor mulr_3_453 xor mulr_4_453;
sumr_454<= mulr_1_454 xor mulr_2_454 xor mulr_3_454 xor mulr_4_454;
sumr_455<= mulr_1_455 xor mulr_2_455 xor mulr_3_455 xor mulr_4_455;
sumr_456<= mulr_1_456 xor mulr_2_456 xor mulr_3_456 xor mulr_4_456;
sumr_457<= mulr_1_457 xor mulr_2_457 xor mulr_3_457 xor mulr_4_457;
sumr_458<= mulr_1_458 xor mulr_2_458 xor mulr_3_458 xor mulr_4_458;
sumr_459<= mulr_1_459 xor mulr_2_459 xor mulr_3_459 xor mulr_4_459;
sumr_460<= mulr_1_460 xor mulr_2_460 xor mulr_3_460 xor mulr_4_460;
sumr_461<= mulr_1_461 xor mulr_2_461 xor mulr_3_461 xor mulr_4_461;
sumr_462<= mulr_1_462 xor mulr_2_462 xor mulr_3_462 xor mulr_4_462;
sumr_463<= mulr_1_463 xor mulr_2_463 xor mulr_3_463 xor mulr_4_463;
sumr_464<= mulr_1_464 xor mulr_2_464 xor mulr_3_464 xor mulr_4_464;
sumr_465<= mulr_1_465 xor mulr_2_465 xor mulr_3_465 xor mulr_4_465;
sumr_466<= mulr_1_466 xor mulr_2_466 xor mulr_3_466 xor mulr_4_466;
sumr_467<= mulr_1_467 xor mulr_2_467 xor mulr_3_467 xor mulr_4_467;
sumr_468<= mulr_1_468 xor mulr_2_468 xor mulr_3_468 xor mulr_4_468;
sumr_469<= mulr_1_469 xor mulr_2_469 xor mulr_3_469 xor mulr_4_469;
sumr_470<= mulr_1_470 xor mulr_2_470 xor mulr_3_470 xor mulr_4_470;
sumr_471<= mulr_1_471 xor mulr_2_471 xor mulr_3_471 xor mulr_4_471;
sumr_472<= mulr_1_472 xor mulr_2_472 xor mulr_3_472 xor mulr_4_472;
sumr_473<= mulr_1_473 xor mulr_2_473 xor mulr_3_473 xor mulr_4_473;
sumr_474<= mulr_1_474 xor mulr_2_474 xor mulr_3_474 xor mulr_4_474;
sumr_475<= mulr_1_475 xor mulr_2_475 xor mulr_3_475 xor mulr_4_475;
sumr_476<= mulr_1_476 xor mulr_2_476 xor mulr_3_476 xor mulr_4_476;
sumr_477<= mulr_1_477 xor mulr_2_477 xor mulr_3_477 xor mulr_4_477;
sumr_478<= mulr_1_478 xor mulr_2_478 xor mulr_3_478 xor mulr_4_478;
sumr_479<= mulr_1_479 xor mulr_2_479 xor mulr_3_479 xor mulr_4_479;
sumr_480<= mulr_1_480 xor mulr_2_480 xor mulr_3_480 xor mulr_4_480;
sumr_481<= mulr_1_481 xor mulr_2_481 xor mulr_3_481 xor mulr_4_481;
sumr_482<= mulr_1_482 xor mulr_2_482 xor mulr_3_482 xor mulr_4_482;
sumr_483<= mulr_1_483 xor mulr_2_483 xor mulr_3_483 xor mulr_4_483;
sumr_484<= mulr_1_484 xor mulr_2_484 xor mulr_3_484 xor mulr_4_484;
sumr_485<= mulr_1_485 xor mulr_2_485 xor mulr_3_485 xor mulr_4_485;
sumr_486<= mulr_1_486 xor mulr_2_486 xor mulr_3_486 xor mulr_4_486;
sumr_487<= mulr_1_487 xor mulr_2_487 xor mulr_3_487 xor mulr_4_487;
sumr_488<= mulr_1_488 xor mulr_2_488 xor mulr_3_488 xor mulr_4_488;
sumr_489<= mulr_1_489 xor mulr_2_489 xor mulr_3_489 xor mulr_4_489;
sumr_490<= mulr_1_490 xor mulr_2_490 xor mulr_3_490 xor mulr_4_490;
sumr_491<= mulr_1_491 xor mulr_2_491 xor mulr_3_491 xor mulr_4_491;
sumr_492<= mulr_1_492 xor mulr_2_492 xor mulr_3_492 xor mulr_4_492;
sumr_493<= mulr_1_493 xor mulr_2_493 xor mulr_3_493 xor mulr_4_493;
sumr_494<= mulr_1_494 xor mulr_2_494 xor mulr_3_494 xor mulr_4_494;
sumr_495<= mulr_1_495 xor mulr_2_495 xor mulr_3_495 xor mulr_4_495;
sumr_496<= mulr_1_496 xor mulr_2_496 xor mulr_3_496 xor mulr_4_496;
sumr_497<= mulr_1_497 xor mulr_2_497 xor mulr_3_497 xor mulr_4_497;
sumr_498<= mulr_1_498 xor mulr_2_498 xor mulr_3_498 xor mulr_4_498;
sumr_499<= mulr_1_499 xor mulr_2_499 xor mulr_3_499 xor mulr_4_499;
sumr_500<= mulr_1_500 xor mulr_2_500 xor mulr_3_500 xor mulr_4_500;
sumr_501<= mulr_1_501 xor mulr_2_501 xor mulr_3_501 xor mulr_4_501;
sumr_502<= mulr_1_502 xor mulr_2_502 xor mulr_3_502 xor mulr_4_502;
sumr_503<= mulr_1_503 xor mulr_2_503 xor mulr_3_503 xor mulr_4_503;
sumr_504<= mulr_1_504 xor mulr_2_504 xor mulr_3_504 xor mulr_4_504;
sumr_505<= mulr_1_505 xor mulr_2_505 xor mulr_3_505 xor mulr_4_505;
sumr_506<= mulr_1_506 xor mulr_2_506 xor mulr_3_506 xor mulr_4_506;
sumr_507<= mulr_1_507 xor mulr_2_507 xor mulr_3_507 xor mulr_4_507;
sumr_508<= mulr_1_508 xor mulr_2_508 xor mulr_3_508 xor mulr_4_508;
sumr_509<= mulr_1_509 xor mulr_2_509 xor mulr_3_509 xor mulr_4_509;
sumr_510<= mulr_1_510 xor mulr_2_510 xor mulr_3_510 xor mulr_4_510;
sumr_511<= mulr_1_511 xor mulr_2_511 xor mulr_3_511 xor mulr_4_511;
sumr_512<= mulr_1_512 xor mulr_2_512 xor mulr_3_512 xor mulr_4_512;
sumr_513<= mulr_1_513 xor mulr_2_513 xor mulr_3_513 xor mulr_4_513;
sumr_514<= mulr_1_514 xor mulr_2_514 xor mulr_3_514 xor mulr_4_514;
sumr_515<= mulr_1_515 xor mulr_2_515 xor mulr_3_515 xor mulr_4_515;
sumr_516<= mulr_1_516 xor mulr_2_516 xor mulr_3_516 xor mulr_4_516;
sumr_517<= mulr_1_517 xor mulr_2_517 xor mulr_3_517 xor mulr_4_517;
sumr_518<= mulr_1_518 xor mulr_2_518 xor mulr_3_518 xor mulr_4_518;
sumr_519<= mulr_1_519 xor mulr_2_519 xor mulr_3_519 xor mulr_4_519;
sumr_520<= mulr_1_520 xor mulr_2_520 xor mulr_3_520 xor mulr_4_520;
sumr_521<= mulr_1_521 xor mulr_2_521 xor mulr_3_521 xor mulr_4_521;
sumr_522<= mulr_1_522 xor mulr_2_522 xor mulr_3_522 xor mulr_4_522;
sumr_523<= mulr_1_523 xor mulr_2_523 xor mulr_3_523 xor mulr_4_523;
sumr_524<= mulr_1_524 xor mulr_2_524 xor mulr_3_524 xor mulr_4_524;
sumr_525<= mulr_1_525 xor mulr_2_525 xor mulr_3_525 xor mulr_4_525;
sumr_526<= mulr_1_526 xor mulr_2_526 xor mulr_3_526 xor mulr_4_526;
sumr_527<= mulr_1_527 xor mulr_2_527 xor mulr_3_527 xor mulr_4_527;
sumr_528<= mulr_1_528 xor mulr_2_528 xor mulr_3_528 xor mulr_4_528;
sumr_529<= mulr_1_529 xor mulr_2_529 xor mulr_3_529 xor mulr_4_529;
sumr_530<= mulr_1_530 xor mulr_2_530 xor mulr_3_530 xor mulr_4_530;
sumr_531<= mulr_1_531 xor mulr_2_531 xor mulr_3_531 xor mulr_4_531;
sumr_532<= mulr_1_532 xor mulr_2_532 xor mulr_3_532 xor mulr_4_532;
sumr_533<= mulr_1_533 xor mulr_2_533 xor mulr_3_533 xor mulr_4_533;
sumr_534<= mulr_1_534 xor mulr_2_534 xor mulr_3_534 xor mulr_4_534;
sumr_535<= mulr_1_535 xor mulr_2_535 xor mulr_3_535 xor mulr_4_535;
sumr_536<= mulr_1_536 xor mulr_2_536 xor mulr_3_536 xor mulr_4_536;
sumr_537<= mulr_1_537 xor mulr_2_537 xor mulr_3_537 xor mulr_4_537;
sumr_538<= mulr_1_538 xor mulr_2_538 xor mulr_3_538 xor mulr_4_538;
sumr_539<= mulr_1_539 xor mulr_2_539 xor mulr_3_539 xor mulr_4_539;
sumr_540<= mulr_1_540 xor mulr_2_540 xor mulr_3_540 xor mulr_4_540;
sumr_541<= mulr_1_541 xor mulr_2_541 xor mulr_3_541 xor mulr_4_541;
sumr_542<= mulr_1_542 xor mulr_2_542 xor mulr_3_542 xor mulr_4_542;
sumr_543<= mulr_1_543 xor mulr_2_543 xor mulr_3_543 xor mulr_4_543;
sumr_544<= mulr_1_544 xor mulr_2_544 xor mulr_3_544 xor mulr_4_544;
sumr_545<= mulr_1_545 xor mulr_2_545 xor mulr_3_545 xor mulr_4_545;
sumr_546<= mulr_1_546 xor mulr_2_546 xor mulr_3_546 xor mulr_4_546;
sumr_547<= mulr_1_547 xor mulr_2_547 xor mulr_3_547 xor mulr_4_547;
sumr_548<= mulr_1_548 xor mulr_2_548 xor mulr_3_548 xor mulr_4_548;
sumr_549<= mulr_1_549 xor mulr_2_549 xor mulr_3_549 xor mulr_4_549;
sumr_550<= mulr_1_550 xor mulr_2_550 xor mulr_3_550 xor mulr_4_550;
sumr_551<= mulr_1_551 xor mulr_2_551 xor mulr_3_551 xor mulr_4_551;
sumr_552<= mulr_1_552 xor mulr_2_552 xor mulr_3_552 xor mulr_4_552;
sumr_553<= mulr_1_553 xor mulr_2_553 xor mulr_3_553 xor mulr_4_553;
sumr_554<= mulr_1_554 xor mulr_2_554 xor mulr_3_554 xor mulr_4_554;
sumr_555<= mulr_1_555 xor mulr_2_555 xor mulr_3_555 xor mulr_4_555;
sumr_556<= mulr_1_556 xor mulr_2_556 xor mulr_3_556 xor mulr_4_556;
sumr_557<= mulr_1_557 xor mulr_2_557 xor mulr_3_557 xor mulr_4_557;
sumr_558<= mulr_1_558 xor mulr_2_558 xor mulr_3_558 xor mulr_4_558;
sumr_559<= mulr_1_559 xor mulr_2_559 xor mulr_3_559 xor mulr_4_559;
sumr_560<= mulr_1_560 xor mulr_2_560 xor mulr_3_560 xor mulr_4_560;
sumr_561<= mulr_1_561 xor mulr_2_561 xor mulr_3_561 xor mulr_4_561;
sumr_562<= mulr_1_562 xor mulr_2_562 xor mulr_3_562 xor mulr_4_562;
sumr_563<= mulr_1_563 xor mulr_2_563 xor mulr_3_563 xor mulr_4_563;
sumr_564<= mulr_1_564 xor mulr_2_564 xor mulr_3_564 xor mulr_4_564;
sumr_565<= mulr_1_565 xor mulr_2_565 xor mulr_3_565 xor mulr_4_565;
sumr_566<= mulr_1_566 xor mulr_2_566 xor mulr_3_566 xor mulr_4_566;
sumr_567<= mulr_1_567 xor mulr_2_567 xor mulr_3_567 xor mulr_4_567;
sumr_568<= mulr_1_568 xor mulr_2_568 xor mulr_3_568 xor mulr_4_568;
sumr_569<= mulr_1_569 xor mulr_2_569 xor mulr_3_569 xor mulr_4_569;
sumr_570<= mulr_1_570 xor mulr_2_570 xor mulr_3_570 xor mulr_4_570;
sumr_571<= mulr_1_571 xor mulr_2_571 xor mulr_3_571 xor mulr_4_571;
sumr_572<= mulr_1_572 xor mulr_2_572 xor mulr_3_572 xor mulr_4_572;
sumr_573<= mulr_1_573 xor mulr_2_573 xor mulr_3_573 xor mulr_4_573;
sumr_574<= mulr_1_574 xor mulr_2_574 xor mulr_3_574 xor mulr_4_574;
sumr_575<= mulr_1_575 xor mulr_2_575 xor mulr_3_575 xor mulr_4_575;
sumr_576<= mulr_1_576 xor mulr_2_576 xor mulr_3_576 xor mulr_4_576;
sumr_577<= mulr_1_577 xor mulr_2_577 xor mulr_3_577 xor mulr_4_577;
sumr_578<= mulr_1_578 xor mulr_2_578 xor mulr_3_578 xor mulr_4_578;
sumr_579<= mulr_1_579 xor mulr_2_579 xor mulr_3_579 xor mulr_4_579;
sumr_580<= mulr_1_580 xor mulr_2_580 xor mulr_3_580 xor mulr_4_580;
sumr_581<= mulr_1_581 xor mulr_2_581 xor mulr_3_581 xor mulr_4_581;
sumr_582<= mulr_1_582 xor mulr_2_582 xor mulr_3_582 xor mulr_4_582;
sumr_583<= mulr_1_583 xor mulr_2_583 xor mulr_3_583 xor mulr_4_583;
sumr_584<= mulr_1_584 xor mulr_2_584 xor mulr_3_584 xor mulr_4_584;
sumr_585<= mulr_1_585 xor mulr_2_585 xor mulr_3_585 xor mulr_4_585;
sumr_586<= mulr_1_586 xor mulr_2_586 xor mulr_3_586 xor mulr_4_586;
sumr_587<= mulr_1_587 xor mulr_2_587 xor mulr_3_587 xor mulr_4_587;
sumr_588<= mulr_1_588 xor mulr_2_588 xor mulr_3_588 xor mulr_4_588;
sumr_589<= mulr_1_589 xor mulr_2_589 xor mulr_3_589 xor mulr_4_589;
sumr_590<= mulr_1_590 xor mulr_2_590 xor mulr_3_590 xor mulr_4_590;
sumr_591<= mulr_1_591 xor mulr_2_591 xor mulr_3_591 xor mulr_4_591;
sumr_592<= mulr_1_592 xor mulr_2_592 xor mulr_3_592 xor mulr_4_592;
sumr_593<= mulr_1_593 xor mulr_2_593 xor mulr_3_593 xor mulr_4_593;
sumr_594<= mulr_1_594 xor mulr_2_594 xor mulr_3_594 xor mulr_4_594;
sumr_595<= mulr_1_595 xor mulr_2_595 xor mulr_3_595 xor mulr_4_595;
sumr_596<= mulr_1_596 xor mulr_2_596 xor mulr_3_596 xor mulr_4_596;
sumr_597<= mulr_1_597 xor mulr_2_597 xor mulr_3_597 xor mulr_4_597;
sumr_598<= mulr_1_598 xor mulr_2_598 xor mulr_3_598 xor mulr_4_598;
sumr_599<= mulr_1_599 xor mulr_2_599 xor mulr_3_599 xor mulr_4_599;
sumr_600<= mulr_1_600 xor mulr_2_600 xor mulr_3_600 xor mulr_4_600;
sumr_601<= mulr_1_601 xor mulr_2_601 xor mulr_3_601 xor mulr_4_601;
sumr_602<= mulr_1_602 xor mulr_2_602 xor mulr_3_602 xor mulr_4_602;
sumr_603<= mulr_1_603 xor mulr_2_603 xor mulr_3_603 xor mulr_4_603;
sumr_604<= mulr_1_604 xor mulr_2_604 xor mulr_3_604 xor mulr_4_604;
sumr_605<= mulr_1_605 xor mulr_2_605 xor mulr_3_605 xor mulr_4_605;
sumr_606<= mulr_1_606 xor mulr_2_606 xor mulr_3_606 xor mulr_4_606;
sumr_607<= mulr_1_607 xor mulr_2_607 xor mulr_3_607 xor mulr_4_607;
sumr_608<= mulr_1_608 xor mulr_2_608 xor mulr_3_608 xor mulr_4_608;
sumr_609<= mulr_1_609 xor mulr_2_609 xor mulr_3_609 xor mulr_4_609;
sumr_610<= mulr_1_610 xor mulr_2_610 xor mulr_3_610 xor mulr_4_610;
sumr_611<= mulr_1_611 xor mulr_2_611 xor mulr_3_611 xor mulr_4_611;
sumr_612<= mulr_1_612 xor mulr_2_612 xor mulr_3_612 xor mulr_4_612;
sumr_613<= mulr_1_613 xor mulr_2_613 xor mulr_3_613 xor mulr_4_613;
sumr_614<= mulr_1_614 xor mulr_2_614 xor mulr_3_614 xor mulr_4_614;
sumr_615<= mulr_1_615 xor mulr_2_615 xor mulr_3_615 xor mulr_4_615;
sumr_616<= mulr_1_616 xor mulr_2_616 xor mulr_3_616 xor mulr_4_616;
sumr_617<= mulr_1_617 xor mulr_2_617 xor mulr_3_617 xor mulr_4_617;
sumr_618<= mulr_1_618 xor mulr_2_618 xor mulr_3_618 xor mulr_4_618;
sumr_619<= mulr_1_619 xor mulr_2_619 xor mulr_3_619 xor mulr_4_619;
sumr_620<= mulr_1_620 xor mulr_2_620 xor mulr_3_620 xor mulr_4_620;
sumr_621<= mulr_1_621 xor mulr_2_621 xor mulr_3_621 xor mulr_4_621;
sumr_622<= mulr_1_622 xor mulr_2_622 xor mulr_3_622 xor mulr_4_622;
sumr_623<= mulr_1_623 xor mulr_2_623 xor mulr_3_623 xor mulr_4_623;
sumr_624<= mulr_1_624 xor mulr_2_624 xor mulr_3_624 xor mulr_4_624;
sumr_625<= mulr_1_625 xor mulr_2_625 xor mulr_3_625 xor mulr_4_625;
sumr_626<= mulr_1_626 xor mulr_2_626 xor mulr_3_626 xor mulr_4_626;
sumr_627<= mulr_1_627 xor mulr_2_627 xor mulr_3_627 xor mulr_4_627;
sumr_628<= mulr_1_628 xor mulr_2_628 xor mulr_3_628 xor mulr_4_628;
sumr_629<= mulr_1_629 xor mulr_2_629 xor mulr_3_629 xor mulr_4_629;
sumr_630<= mulr_1_630 xor mulr_2_630 xor mulr_3_630 xor mulr_4_630;
sumr_631<= mulr_1_631 xor mulr_2_631 xor mulr_3_631 xor mulr_4_631;
sumr_632<= mulr_1_632 xor mulr_2_632 xor mulr_3_632 xor mulr_4_632;
sumr_633<= mulr_1_633 xor mulr_2_633 xor mulr_3_633 xor mulr_4_633;
sumr_634<= mulr_1_634 xor mulr_2_634 xor mulr_3_634 xor mulr_4_634;
sumr_635<= mulr_1_635 xor mulr_2_635 xor mulr_3_635 xor mulr_4_635;
sumr_636<= mulr_1_636 xor mulr_2_636 xor mulr_3_636 xor mulr_4_636;
sumr_637<= mulr_1_637 xor mulr_2_637 xor mulr_3_637 xor mulr_4_637;
sumr_638<= mulr_1_638 xor mulr_2_638 xor mulr_3_638 xor mulr_4_638;
sumr_639<= mulr_1_639 xor mulr_2_639 xor mulr_3_639 xor mulr_4_639;
sumr_640<= mulr_1_640 xor mulr_2_640 xor mulr_3_640 xor mulr_4_640;
sumr_641<= mulr_1_641 xor mulr_2_641 xor mulr_3_641 xor mulr_4_641;
sumr_642<= mulr_1_642 xor mulr_2_642 xor mulr_3_642 xor mulr_4_642;
sumr_643<= mulr_1_643 xor mulr_2_643 xor mulr_3_643 xor mulr_4_643;
sumr_644<= mulr_1_644 xor mulr_2_644 xor mulr_3_644 xor mulr_4_644;
sumr_645<= mulr_1_645 xor mulr_2_645 xor mulr_3_645 xor mulr_4_645;
sumr_646<= mulr_1_646 xor mulr_2_646 xor mulr_3_646 xor mulr_4_646;
sumr_647<= mulr_1_647 xor mulr_2_647 xor mulr_3_647 xor mulr_4_647;
sumr_648<= mulr_1_648 xor mulr_2_648 xor mulr_3_648 xor mulr_4_648;
sumr_649<= mulr_1_649 xor mulr_2_649 xor mulr_3_649 xor mulr_4_649;
sumr_650<= mulr_1_650 xor mulr_2_650 xor mulr_3_650 xor mulr_4_650;
sumr_651<= mulr_1_651 xor mulr_2_651 xor mulr_3_651 xor mulr_4_651;
sumr_652<= mulr_1_652 xor mulr_2_652 xor mulr_3_652 xor mulr_4_652;
sumr_653<= mulr_1_653 xor mulr_2_653 xor mulr_3_653 xor mulr_4_653;
sumr_654<= mulr_1_654 xor mulr_2_654 xor mulr_3_654 xor mulr_4_654;
sumr_655<= mulr_1_655 xor mulr_2_655 xor mulr_3_655 xor mulr_4_655;
sumr_656<= mulr_1_656 xor mulr_2_656 xor mulr_3_656 xor mulr_4_656;
sumr_657<= mulr_1_657 xor mulr_2_657 xor mulr_3_657 xor mulr_4_657;
sumr_658<= mulr_1_658 xor mulr_2_658 xor mulr_3_658 xor mulr_4_658;
sumr_659<= mulr_1_659 xor mulr_2_659 xor mulr_3_659 xor mulr_4_659;
sumr_660<= mulr_1_660 xor mulr_2_660 xor mulr_3_660 xor mulr_4_660;
sumr_661<= mulr_1_661 xor mulr_2_661 xor mulr_3_661 xor mulr_4_661;
sumr_662<= mulr_1_662 xor mulr_2_662 xor mulr_3_662 xor mulr_4_662;
sumr_663<= mulr_1_663 xor mulr_2_663 xor mulr_3_663 xor mulr_4_663;
sumr_664<= mulr_1_664 xor mulr_2_664 xor mulr_3_664 xor mulr_4_664;
sumr_665<= mulr_1_665 xor mulr_2_665 xor mulr_3_665 xor mulr_4_665;
sumr_666<= mulr_1_666 xor mulr_2_666 xor mulr_3_666 xor mulr_4_666;
sumr_667<= mulr_1_667 xor mulr_2_667 xor mulr_3_667 xor mulr_4_667;
sumr_668<= mulr_1_668 xor mulr_2_668 xor mulr_3_668 xor mulr_4_668;
sumr_669<= mulr_1_669 xor mulr_2_669 xor mulr_3_669 xor mulr_4_669;
sumr_670<= mulr_1_670 xor mulr_2_670 xor mulr_3_670 xor mulr_4_670;
sumr_671<= mulr_1_671 xor mulr_2_671 xor mulr_3_671 xor mulr_4_671;
sumr_672<= mulr_1_672 xor mulr_2_672 xor mulr_3_672 xor mulr_4_672;
sumr_673<= mulr_1_673 xor mulr_2_673 xor mulr_3_673 xor mulr_4_673;
sumr_674<= mulr_1_674 xor mulr_2_674 xor mulr_3_674 xor mulr_4_674;
sumr_675<= mulr_1_675 xor mulr_2_675 xor mulr_3_675 xor mulr_4_675;
sumr_676<= mulr_1_676 xor mulr_2_676 xor mulr_3_676 xor mulr_4_676;
sumr_677<= mulr_1_677 xor mulr_2_677 xor mulr_3_677 xor mulr_4_677;
sumr_678<= mulr_1_678 xor mulr_2_678 xor mulr_3_678 xor mulr_4_678;
sumr_679<= mulr_1_679 xor mulr_2_679 xor mulr_3_679 xor mulr_4_679;
sumr_680<= mulr_1_680 xor mulr_2_680 xor mulr_3_680 xor mulr_4_680;
sumr_681<= mulr_1_681 xor mulr_2_681 xor mulr_3_681 xor mulr_4_681;
sumr_682<= mulr_1_682 xor mulr_2_682 xor mulr_3_682 xor mulr_4_682;
sumr_683<= mulr_1_683 xor mulr_2_683 xor mulr_3_683 xor mulr_4_683;
sumr_684<= mulr_1_684 xor mulr_2_684 xor mulr_3_684 xor mulr_4_684;
sumr_685<= mulr_1_685 xor mulr_2_685 xor mulr_3_685 xor mulr_4_685;
sumr_686<= mulr_1_686 xor mulr_2_686 xor mulr_3_686 xor mulr_4_686;
sumr_687<= mulr_1_687 xor mulr_2_687 xor mulr_3_687 xor mulr_4_687;
sumr_688<= mulr_1_688 xor mulr_2_688 xor mulr_3_688 xor mulr_4_688;
sumr_689<= mulr_1_689 xor mulr_2_689 xor mulr_3_689 xor mulr_4_689;
sumr_690<= mulr_1_690 xor mulr_2_690 xor mulr_3_690 xor mulr_4_690;
sumr_691<= mulr_1_691 xor mulr_2_691 xor mulr_3_691 xor mulr_4_691;
sumr_692<= mulr_1_692 xor mulr_2_692 xor mulr_3_692 xor mulr_4_692;
sumr_693<= mulr_1_693 xor mulr_2_693 xor mulr_3_693 xor mulr_4_693;
sumr_694<= mulr_1_694 xor mulr_2_694 xor mulr_3_694 xor mulr_4_694;
sumr_695<= mulr_1_695 xor mulr_2_695 xor mulr_3_695 xor mulr_4_695;
sumr_696<= mulr_1_696 xor mulr_2_696 xor mulr_3_696 xor mulr_4_696;
sumr_697<= mulr_1_697 xor mulr_2_697 xor mulr_3_697 xor mulr_4_697;
sumr_698<= mulr_1_698 xor mulr_2_698 xor mulr_3_698 xor mulr_4_698;
sumr_699<= mulr_1_699 xor mulr_2_699 xor mulr_3_699 xor mulr_4_699;
sumr_700<= mulr_1_700 xor mulr_2_700 xor mulr_3_700 xor mulr_4_700;
sumr_701<= mulr_1_701 xor mulr_2_701 xor mulr_3_701 xor mulr_4_701;
sumr_702<= mulr_1_702 xor mulr_2_702 xor mulr_3_702 xor mulr_4_702;
sumr_703<= mulr_1_703 xor mulr_2_703 xor mulr_3_703 xor mulr_4_703;
sumr_704<= mulr_1_704 xor mulr_2_704 xor mulr_3_704 xor mulr_4_704;
sumr_705<= mulr_1_705 xor mulr_2_705 xor mulr_3_705 xor mulr_4_705;
sumr_706<= mulr_1_706 xor mulr_2_706 xor mulr_3_706 xor mulr_4_706;
sumr_707<= mulr_1_707 xor mulr_2_707 xor mulr_3_707 xor mulr_4_707;
sumr_708<= mulr_1_708 xor mulr_2_708 xor mulr_3_708 xor mulr_4_708;
sumr_709<= mulr_1_709 xor mulr_2_709 xor mulr_3_709 xor mulr_4_709;
sumr_710<= mulr_1_710 xor mulr_2_710 xor mulr_3_710 xor mulr_4_710;
sumr_711<= mulr_1_711 xor mulr_2_711 xor mulr_3_711 xor mulr_4_711;
sumr_712<= mulr_1_712 xor mulr_2_712 xor mulr_3_712 xor mulr_4_712;
sumr_713<= mulr_1_713 xor mulr_2_713 xor mulr_3_713 xor mulr_4_713;
sumr_714<= mulr_1_714 xor mulr_2_714 xor mulr_3_714 xor mulr_4_714;
sumr_715<= mulr_1_715 xor mulr_2_715 xor mulr_3_715 xor mulr_4_715;
sumr_716<= mulr_1_716 xor mulr_2_716 xor mulr_3_716 xor mulr_4_716;
sumr_717<= mulr_1_717 xor mulr_2_717 xor mulr_3_717 xor mulr_4_717;
sumr_718<= mulr_1_718 xor mulr_2_718 xor mulr_3_718 xor mulr_4_718;
sumr_719<= mulr_1_719 xor mulr_2_719 xor mulr_3_719 xor mulr_4_719;
sumr_720<= mulr_1_720 xor mulr_2_720 xor mulr_3_720 xor mulr_4_720;
sumr_721<= mulr_1_721 xor mulr_2_721 xor mulr_3_721 xor mulr_4_721;
sumr_722<= mulr_1_722 xor mulr_2_722 xor mulr_3_722 xor mulr_4_722;
sumr_723<= mulr_1_723 xor mulr_2_723 xor mulr_3_723 xor mulr_4_723;
sumr_724<= mulr_1_724 xor mulr_2_724 xor mulr_3_724 xor mulr_4_724;
sumr_725<= mulr_1_725 xor mulr_2_725 xor mulr_3_725 xor mulr_4_725;
sumr_726<= mulr_1_726 xor mulr_2_726 xor mulr_3_726 xor mulr_4_726;
sumr_727<= mulr_1_727 xor mulr_2_727 xor mulr_3_727 xor mulr_4_727;
sumr_728<= mulr_1_728 xor mulr_2_728 xor mulr_3_728 xor mulr_4_728;
sumr_729<= mulr_1_729 xor mulr_2_729 xor mulr_3_729 xor mulr_4_729;
sumr_730<= mulr_1_730 xor mulr_2_730 xor mulr_3_730 xor mulr_4_730;
sumr_731<= mulr_1_731 xor mulr_2_731 xor mulr_3_731 xor mulr_4_731;
sumr_732<= mulr_1_732 xor mulr_2_732 xor mulr_3_732 xor mulr_4_732;
sumr_733<= mulr_1_733 xor mulr_2_733 xor mulr_3_733 xor mulr_4_733;
sumr_734<= mulr_1_734 xor mulr_2_734 xor mulr_3_734 xor mulr_4_734;
sumr_735<= mulr_1_735 xor mulr_2_735 xor mulr_3_735 xor mulr_4_735;
sumr_736<= mulr_1_736 xor mulr_2_736 xor mulr_3_736 xor mulr_4_736;
sumr_737<= mulr_1_737 xor mulr_2_737 xor mulr_3_737 xor mulr_4_737;
sumr_738<= mulr_1_738 xor mulr_2_738 xor mulr_3_738 xor mulr_4_738;
sumr_739<= mulr_1_739 xor mulr_2_739 xor mulr_3_739 xor mulr_4_739;
sumr_740<= mulr_1_740 xor mulr_2_740 xor mulr_3_740 xor mulr_4_740;
sumr_741<= mulr_1_741 xor mulr_2_741 xor mulr_3_741 xor mulr_4_741;
sumr_742<= mulr_1_742 xor mulr_2_742 xor mulr_3_742 xor mulr_4_742;
sumr_743<= mulr_1_743 xor mulr_2_743 xor mulr_3_743 xor mulr_4_743;
sumr_744<= mulr_1_744 xor mulr_2_744 xor mulr_3_744 xor mulr_4_744;
sumr_745<= mulr_1_745 xor mulr_2_745 xor mulr_3_745 xor mulr_4_745;
sumr_746<= mulr_1_746 xor mulr_2_746 xor mulr_3_746 xor mulr_4_746;
sumr_747<= mulr_1_747 xor mulr_2_747 xor mulr_3_747 xor mulr_4_747;
sumr_748<= mulr_1_748 xor mulr_2_748 xor mulr_3_748 xor mulr_4_748;
sumr_749<= mulr_1_749 xor mulr_2_749 xor mulr_3_749 xor mulr_4_749;
sumr_750<= mulr_1_750 xor mulr_2_750 xor mulr_3_750 xor mulr_4_750;
sumr_751<= mulr_1_751 xor mulr_2_751 xor mulr_3_751 xor mulr_4_751;
sumr_752<= mulr_1_752 xor mulr_2_752 xor mulr_3_752 xor mulr_4_752;
sumr_753<= mulr_1_753 xor mulr_2_753 xor mulr_3_753 xor mulr_4_753;
sumr_754<= mulr_1_754 xor mulr_2_754 xor mulr_3_754 xor mulr_4_754;
sumr_755<= mulr_1_755 xor mulr_2_755 xor mulr_3_755 xor mulr_4_755;
sumr_756<= mulr_1_756 xor mulr_2_756 xor mulr_3_756 xor mulr_4_756;
sumr_757<= mulr_1_757 xor mulr_2_757 xor mulr_3_757 xor mulr_4_757;
sumr_758<= mulr_1_758 xor mulr_2_758 xor mulr_3_758 xor mulr_4_758;
sumr_759<= mulr_1_759 xor mulr_2_759 xor mulr_3_759 xor mulr_4_759;
sumr_760<= mulr_1_760 xor mulr_2_760 xor mulr_3_760 xor mulr_4_760;
sumr_761<= mulr_1_761 xor mulr_2_761 xor mulr_3_761 xor mulr_4_761;
sumr_762<= mulr_1_762 xor mulr_2_762 xor mulr_3_762 xor mulr_4_762;
sumr_763<= mulr_1_763 xor mulr_2_763 xor mulr_3_763 xor mulr_4_763;
sumr_764<= mulr_1_764 xor mulr_2_764 xor mulr_3_764 xor mulr_4_764;
sumr_765<= mulr_1_765 xor mulr_2_765 xor mulr_3_765 xor mulr_4_765;
sumr_766<= mulr_1_766 xor mulr_2_766 xor mulr_3_766 xor mulr_4_766;
sumr_767<= mulr_1_767 xor mulr_2_767 xor mulr_3_767 xor mulr_4_767;
sumr_768<= mulr_1_768 xor mulr_2_768 xor mulr_3_768 xor mulr_4_768;
sumr_769<= mulr_1_769 xor mulr_2_769 xor mulr_3_769 xor mulr_4_769;
sumr_770<= mulr_1_770 xor mulr_2_770 xor mulr_3_770 xor mulr_4_770;
sumr_771<= mulr_1_771 xor mulr_2_771 xor mulr_3_771 xor mulr_4_771;
sumr_772<= mulr_1_772 xor mulr_2_772 xor mulr_3_772 xor mulr_4_772;
sumr_773<= mulr_1_773 xor mulr_2_773 xor mulr_3_773 xor mulr_4_773;
sumr_774<= mulr_1_774 xor mulr_2_774 xor mulr_3_774 xor mulr_4_774;
sumr_775<= mulr_1_775 xor mulr_2_775 xor mulr_3_775 xor mulr_4_775;
sumr_776<= mulr_1_776 xor mulr_2_776 xor mulr_3_776 xor mulr_4_776;
sumr_777<= mulr_1_777 xor mulr_2_777 xor mulr_3_777 xor mulr_4_777;
sumr_778<= mulr_1_778 xor mulr_2_778 xor mulr_3_778 xor mulr_4_778;
sumr_779<= mulr_1_779 xor mulr_2_779 xor mulr_3_779 xor mulr_4_779;
sumr_780<= mulr_1_780 xor mulr_2_780 xor mulr_3_780 xor mulr_4_780;
sumr_781<= mulr_1_781 xor mulr_2_781 xor mulr_3_781 xor mulr_4_781;
sumr_782<= mulr_1_782 xor mulr_2_782 xor mulr_3_782 xor mulr_4_782;
sumr_783<= mulr_1_783 xor mulr_2_783 xor mulr_3_783 xor mulr_4_783;
sumr_784<= mulr_1_784 xor mulr_2_784 xor mulr_3_784 xor mulr_4_784;
sumr_785<= mulr_1_785 xor mulr_2_785 xor mulr_3_785 xor mulr_4_785;
sumr_786<= mulr_1_786 xor mulr_2_786 xor mulr_3_786 xor mulr_4_786;
sumr_787<= mulr_1_787 xor mulr_2_787 xor mulr_3_787 xor mulr_4_787;
sumr_788<= mulr_1_788 xor mulr_2_788 xor mulr_3_788 xor mulr_4_788;
sumr_789<= mulr_1_789 xor mulr_2_789 xor mulr_3_789 xor mulr_4_789;
sumr_790<= mulr_1_790 xor mulr_2_790 xor mulr_3_790 xor mulr_4_790;
sumr_791<= mulr_1_791 xor mulr_2_791 xor mulr_3_791 xor mulr_4_791;
sumr_792<= mulr_1_792 xor mulr_2_792 xor mulr_3_792 xor mulr_4_792;
sumr_793<= mulr_1_793 xor mulr_2_793 xor mulr_3_793 xor mulr_4_793;
sumr_794<= mulr_1_794 xor mulr_2_794 xor mulr_3_794 xor mulr_4_794;
sumr_795<= mulr_1_795 xor mulr_2_795 xor mulr_3_795 xor mulr_4_795;
sumr_796<= mulr_1_796 xor mulr_2_796 xor mulr_3_796 xor mulr_4_796;
sumr_797<= mulr_1_797 xor mulr_2_797 xor mulr_3_797 xor mulr_4_797;
sumr_798<= mulr_1_798 xor mulr_2_798 xor mulr_3_798 xor mulr_4_798;
sumr_799<= mulr_1_799 xor mulr_2_799 xor mulr_3_799 xor mulr_4_799;
sumr_800<= mulr_1_800 xor mulr_2_800 xor mulr_3_800 xor mulr_4_800;
sumr_801<= mulr_1_801 xor mulr_2_801 xor mulr_3_801 xor mulr_4_801;
sumr_802<= mulr_1_802 xor mulr_2_802 xor mulr_3_802 xor mulr_4_802;
sumr_803<= mulr_1_803 xor mulr_2_803 xor mulr_3_803 xor mulr_4_803;
sumr_804<= mulr_1_804 xor mulr_2_804 xor mulr_3_804 xor mulr_4_804;
sumr_805<= mulr_1_805 xor mulr_2_805 xor mulr_3_805 xor mulr_4_805;
sumr_806<= mulr_1_806 xor mulr_2_806 xor mulr_3_806 xor mulr_4_806;
sumr_807<= mulr_1_807 xor mulr_2_807 xor mulr_3_807 xor mulr_4_807;
sumr_808<= mulr_1_808 xor mulr_2_808 xor mulr_3_808 xor mulr_4_808;
sumr_809<= mulr_1_809 xor mulr_2_809 xor mulr_3_809 xor mulr_4_809;
sumr_810<= mulr_1_810 xor mulr_2_810 xor mulr_3_810 xor mulr_4_810;
sumr_811<= mulr_1_811 xor mulr_2_811 xor mulr_3_811 xor mulr_4_811;
sumr_812<= mulr_1_812 xor mulr_2_812 xor mulr_3_812 xor mulr_4_812;
sumr_813<= mulr_1_813 xor mulr_2_813 xor mulr_3_813 xor mulr_4_813;
sumr_814<= mulr_1_814 xor mulr_2_814 xor mulr_3_814 xor mulr_4_814;
sumr_815<= mulr_1_815 xor mulr_2_815 xor mulr_3_815 xor mulr_4_815;
sumr_816<= mulr_1_816 xor mulr_2_816 xor mulr_3_816 xor mulr_4_816;
sumr_817<= mulr_1_817 xor mulr_2_817 xor mulr_3_817 xor mulr_4_817;
sumr_818<= mulr_1_818 xor mulr_2_818 xor mulr_3_818 xor mulr_4_818;
sumr_819<= mulr_1_819 xor mulr_2_819 xor mulr_3_819 xor mulr_4_819;
sumr_820<= mulr_1_820 xor mulr_2_820 xor mulr_3_820 xor mulr_4_820;
sumr_821<= mulr_1_821 xor mulr_2_821 xor mulr_3_821 xor mulr_4_821;
sumr_822<= mulr_1_822 xor mulr_2_822 xor mulr_3_822 xor mulr_4_822;
sumr_823<= mulr_1_823 xor mulr_2_823 xor mulr_3_823 xor mulr_4_823;
sumr_824<= mulr_1_824 xor mulr_2_824 xor mulr_3_824 xor mulr_4_824;
sumr_825<= mulr_1_825 xor mulr_2_825 xor mulr_3_825 xor mulr_4_825;
sumr_826<= mulr_1_826 xor mulr_2_826 xor mulr_3_826 xor mulr_4_826;
sumr_827<= mulr_1_827 xor mulr_2_827 xor mulr_3_827 xor mulr_4_827;
sumr_828<= mulr_1_828 xor mulr_2_828 xor mulr_3_828 xor mulr_4_828;
sumr_829<= mulr_1_829 xor mulr_2_829 xor mulr_3_829 xor mulr_4_829;
sumr_830<= mulr_1_830 xor mulr_2_830 xor mulr_3_830 xor mulr_4_830;
sumr_831<= mulr_1_831 xor mulr_2_831 xor mulr_3_831 xor mulr_4_831;
sumr_832<= mulr_1_832 xor mulr_2_832 xor mulr_3_832 xor mulr_4_832;
sumr_833<= mulr_1_833 xor mulr_2_833 xor mulr_3_833 xor mulr_4_833;
sumr_834<= mulr_1_834 xor mulr_2_834 xor mulr_3_834 xor mulr_4_834;
sumr_835<= mulr_1_835 xor mulr_2_835 xor mulr_3_835 xor mulr_4_835;
sumr_836<= mulr_1_836 xor mulr_2_836 xor mulr_3_836 xor mulr_4_836;
sumr_837<= mulr_1_837 xor mulr_2_837 xor mulr_3_837 xor mulr_4_837;
sumr_838<= mulr_1_838 xor mulr_2_838 xor mulr_3_838 xor mulr_4_838;
sumr_839<= mulr_1_839 xor mulr_2_839 xor mulr_3_839 xor mulr_4_839;
sumr_840<= mulr_1_840 xor mulr_2_840 xor mulr_3_840 xor mulr_4_840;
sumr_841<= mulr_1_841 xor mulr_2_841 xor mulr_3_841 xor mulr_4_841;
sumr_842<= mulr_1_842 xor mulr_2_842 xor mulr_3_842 xor mulr_4_842;
sumr_843<= mulr_1_843 xor mulr_2_843 xor mulr_3_843 xor mulr_4_843;
sumr_844<= mulr_1_844 xor mulr_2_844 xor mulr_3_844 xor mulr_4_844;
sumr_845<= mulr_1_845 xor mulr_2_845 xor mulr_3_845 xor mulr_4_845;
sumr_846<= mulr_1_846 xor mulr_2_846 xor mulr_3_846 xor mulr_4_846;
sumr_847<= mulr_1_847 xor mulr_2_847 xor mulr_3_847 xor mulr_4_847;
sumr_848<= mulr_1_848 xor mulr_2_848 xor mulr_3_848 xor mulr_4_848;
sumr_849<= mulr_1_849 xor mulr_2_849 xor mulr_3_849 xor mulr_4_849;
sumr_850<= mulr_1_850 xor mulr_2_850 xor mulr_3_850 xor mulr_4_850;
sumr_851<= mulr_1_851 xor mulr_2_851 xor mulr_3_851 xor mulr_4_851;
sumr_852<= mulr_1_852 xor mulr_2_852 xor mulr_3_852 xor mulr_4_852;
sumr_853<= mulr_1_853 xor mulr_2_853 xor mulr_3_853 xor mulr_4_853;
sumr_854<= mulr_1_854 xor mulr_2_854 xor mulr_3_854 xor mulr_4_854;
sumr_855<= mulr_1_855 xor mulr_2_855 xor mulr_3_855 xor mulr_4_855;
sumr_856<= mulr_1_856 xor mulr_2_856 xor mulr_3_856 xor mulr_4_856;
sumr_857<= mulr_1_857 xor mulr_2_857 xor mulr_3_857 xor mulr_4_857;
sumr_858<= mulr_1_858 xor mulr_2_858 xor mulr_3_858 xor mulr_4_858;
sumr_859<= mulr_1_859 xor mulr_2_859 xor mulr_3_859 xor mulr_4_859;
sumr_860<= mulr_1_860 xor mulr_2_860 xor mulr_3_860 xor mulr_4_860;
sumr_861<= mulr_1_861 xor mulr_2_861 xor mulr_3_861 xor mulr_4_861;
sumr_862<= mulr_1_862 xor mulr_2_862 xor mulr_3_862 xor mulr_4_862;
sumr_863<= mulr_1_863 xor mulr_2_863 xor mulr_3_863 xor mulr_4_863;
sumr_864<= mulr_1_864 xor mulr_2_864 xor mulr_3_864 xor mulr_4_864;
sumr_865<= mulr_1_865 xor mulr_2_865 xor mulr_3_865 xor mulr_4_865;
sumr_866<= mulr_1_866 xor mulr_2_866 xor mulr_3_866 xor mulr_4_866;
sumr_867<= mulr_1_867 xor mulr_2_867 xor mulr_3_867 xor mulr_4_867;
sumr_868<= mulr_1_868 xor mulr_2_868 xor mulr_3_868 xor mulr_4_868;
sumr_869<= mulr_1_869 xor mulr_2_869 xor mulr_3_869 xor mulr_4_869;
sumr_870<= mulr_1_870 xor mulr_2_870 xor mulr_3_870 xor mulr_4_870;
sumr_871<= mulr_1_871 xor mulr_2_871 xor mulr_3_871 xor mulr_4_871;
sumr_872<= mulr_1_872 xor mulr_2_872 xor mulr_3_872 xor mulr_4_872;
sumr_873<= mulr_1_873 xor mulr_2_873 xor mulr_3_873 xor mulr_4_873;
sumr_874<= mulr_1_874 xor mulr_2_874 xor mulr_3_874 xor mulr_4_874;
sumr_875<= mulr_1_875 xor mulr_2_875 xor mulr_3_875 xor mulr_4_875;
sumr_876<= mulr_1_876 xor mulr_2_876 xor mulr_3_876 xor mulr_4_876;
sumr_877<= mulr_1_877 xor mulr_2_877 xor mulr_3_877 xor mulr_4_877;
sumr_878<= mulr_1_878 xor mulr_2_878 xor mulr_3_878 xor mulr_4_878;
sumr_879<= mulr_1_879 xor mulr_2_879 xor mulr_3_879 xor mulr_4_879;
sumr_880<= mulr_1_880 xor mulr_2_880 xor mulr_3_880 xor mulr_4_880;
sumr_881<= mulr_1_881 xor mulr_2_881 xor mulr_3_881 xor mulr_4_881;
sumr_882<= mulr_1_882 xor mulr_2_882 xor mulr_3_882 xor mulr_4_882;
sumr_883<= mulr_1_883 xor mulr_2_883 xor mulr_3_883 xor mulr_4_883;
sumr_884<= mulr_1_884 xor mulr_2_884 xor mulr_3_884 xor mulr_4_884;
sumr_885<= mulr_1_885 xor mulr_2_885 xor mulr_3_885 xor mulr_4_885;
sumr_886<= mulr_1_886 xor mulr_2_886 xor mulr_3_886 xor mulr_4_886;
sumr_887<= mulr_1_887 xor mulr_2_887 xor mulr_3_887 xor mulr_4_887;
sumr_888<= mulr_1_888 xor mulr_2_888 xor mulr_3_888 xor mulr_4_888;
sumr_889<= mulr_1_889 xor mulr_2_889 xor mulr_3_889 xor mulr_4_889;
sumr_890<= mulr_1_890 xor mulr_2_890 xor mulr_3_890 xor mulr_4_890;
sumr_891<= mulr_1_891 xor mulr_2_891 xor mulr_3_891 xor mulr_4_891;
sumr_892<= mulr_1_892 xor mulr_2_892 xor mulr_3_892 xor mulr_4_892;
sumr_893<= mulr_1_893 xor mulr_2_893 xor mulr_3_893 xor mulr_4_893;
sumr_894<= mulr_1_894 xor mulr_2_894 xor mulr_3_894 xor mulr_4_894;
sumr_895<= mulr_1_895 xor mulr_2_895 xor mulr_3_895 xor mulr_4_895;
sumr_896<= mulr_1_896 xor mulr_2_896 xor mulr_3_896 xor mulr_4_896;
sumr_897<= mulr_1_897 xor mulr_2_897 xor mulr_3_897 xor mulr_4_897;
sumr_898<= mulr_1_898 xor mulr_2_898 xor mulr_3_898 xor mulr_4_898;
sumr_899<= mulr_1_899 xor mulr_2_899 xor mulr_3_899 xor mulr_4_899;
sumr_900<= mulr_1_900 xor mulr_2_900 xor mulr_3_900 xor mulr_4_900;
sumr_901<= mulr_1_901 xor mulr_2_901 xor mulr_3_901 xor mulr_4_901;
sumr_902<= mulr_1_902 xor mulr_2_902 xor mulr_3_902 xor mulr_4_902;
sumr_903<= mulr_1_903 xor mulr_2_903 xor mulr_3_903 xor mulr_4_903;
sumr_904<= mulr_1_904 xor mulr_2_904 xor mulr_3_904 xor mulr_4_904;
sumr_905<= mulr_1_905 xor mulr_2_905 xor mulr_3_905 xor mulr_4_905;
sumr_906<= mulr_1_906 xor mulr_2_906 xor mulr_3_906 xor mulr_4_906;
sumr_907<= mulr_1_907 xor mulr_2_907 xor mulr_3_907 xor mulr_4_907;
sumr_908<= mulr_1_908 xor mulr_2_908 xor mulr_3_908 xor mulr_4_908;
sumr_909<= mulr_1_909 xor mulr_2_909 xor mulr_3_909 xor mulr_4_909;
sumr_910<= mulr_1_910 xor mulr_2_910 xor mulr_3_910 xor mulr_4_910;
sumr_911<= mulr_1_911 xor mulr_2_911 xor mulr_3_911 xor mulr_4_911;
sumr_912<= mulr_1_912 xor mulr_2_912 xor mulr_3_912 xor mulr_4_912;
sumr_913<= mulr_1_913 xor mulr_2_913 xor mulr_3_913 xor mulr_4_913;
sumr_914<= mulr_1_914 xor mulr_2_914 xor mulr_3_914 xor mulr_4_914;
sumr_915<= mulr_1_915 xor mulr_2_915 xor mulr_3_915 xor mulr_4_915;
sumr_916<= mulr_1_916 xor mulr_2_916 xor mulr_3_916 xor mulr_4_916;
sumr_917<= mulr_1_917 xor mulr_2_917 xor mulr_3_917 xor mulr_4_917;
sumr_918<= mulr_1_918 xor mulr_2_918 xor mulr_3_918 xor mulr_4_918;
sumr_919<= mulr_1_919 xor mulr_2_919 xor mulr_3_919 xor mulr_4_919;
sumr_920<= mulr_1_920 xor mulr_2_920 xor mulr_3_920 xor mulr_4_920;
sumr_921<= mulr_1_921 xor mulr_2_921 xor mulr_3_921 xor mulr_4_921;
sumr_922<= mulr_1_922 xor mulr_2_922 xor mulr_3_922 xor mulr_4_922;
sumr_923<= mulr_1_923 xor mulr_2_923 xor mulr_3_923 xor mulr_4_923;
sumr_924<= mulr_1_924 xor mulr_2_924 xor mulr_3_924 xor mulr_4_924;
sumr_925<= mulr_1_925 xor mulr_2_925 xor mulr_3_925 xor mulr_4_925;
sumr_926<= mulr_1_926 xor mulr_2_926 xor mulr_3_926 xor mulr_4_926;
sumr_927<= mulr_1_927 xor mulr_2_927 xor mulr_3_927 xor mulr_4_927;
sumr_928<= mulr_1_928 xor mulr_2_928 xor mulr_3_928 xor mulr_4_928;
sumr_929<= mulr_1_929 xor mulr_2_929 xor mulr_3_929 xor mulr_4_929;
sumr_930<= mulr_1_930 xor mulr_2_930 xor mulr_3_930 xor mulr_4_930;
sumr_931<= mulr_1_931 xor mulr_2_931 xor mulr_3_931 xor mulr_4_931;
sumr_932<= mulr_1_932 xor mulr_2_932 xor mulr_3_932 xor mulr_4_932;
sumr_933<= mulr_1_933 xor mulr_2_933 xor mulr_3_933 xor mulr_4_933;
sumr_934<= mulr_1_934 xor mulr_2_934 xor mulr_3_934 xor mulr_4_934;
sumr_935<= mulr_1_935 xor mulr_2_935 xor mulr_3_935 xor mulr_4_935;
sumr_936<= mulr_1_936 xor mulr_2_936 xor mulr_3_936 xor mulr_4_936;
sumr_937<= mulr_1_937 xor mulr_2_937 xor mulr_3_937 xor mulr_4_937;
sumr_938<= mulr_1_938 xor mulr_2_938 xor mulr_3_938 xor mulr_4_938;
sumr_939<= mulr_1_939 xor mulr_2_939 xor mulr_3_939 xor mulr_4_939;
sumr_940<= mulr_1_940 xor mulr_2_940 xor mulr_3_940 xor mulr_4_940;
sumr_941<= mulr_1_941 xor mulr_2_941 xor mulr_3_941 xor mulr_4_941;
sumr_942<= mulr_1_942 xor mulr_2_942 xor mulr_3_942 xor mulr_4_942;
sumr_943<= mulr_1_943 xor mulr_2_943 xor mulr_3_943 xor mulr_4_943;
sumr_944<= mulr_1_944 xor mulr_2_944 xor mulr_3_944 xor mulr_4_944;
sumr_945<= mulr_1_945 xor mulr_2_945 xor mulr_3_945 xor mulr_4_945;
sumr_946<= mulr_1_946 xor mulr_2_946 xor mulr_3_946 xor mulr_4_946;
sumr_947<= mulr_1_947 xor mulr_2_947 xor mulr_3_947 xor mulr_4_947;
sumr_948<= mulr_1_948 xor mulr_2_948 xor mulr_3_948 xor mulr_4_948;
sumr_949<= mulr_1_949 xor mulr_2_949 xor mulr_3_949 xor mulr_4_949;
sumr_950<= mulr_1_950 xor mulr_2_950 xor mulr_3_950 xor mulr_4_950;
sumr_951<= mulr_1_951 xor mulr_2_951 xor mulr_3_951 xor mulr_4_951;
sumr_952<= mulr_1_952 xor mulr_2_952 xor mulr_3_952 xor mulr_4_952;
sumr_953<= mulr_1_953 xor mulr_2_953 xor mulr_3_953 xor mulr_4_953;
sumr_954<= mulr_1_954 xor mulr_2_954 xor mulr_3_954 xor mulr_4_954;
sumr_955<= mulr_1_955 xor mulr_2_955 xor mulr_3_955 xor mulr_4_955;
sumr_956<= mulr_1_956 xor mulr_2_956 xor mulr_3_956 xor mulr_4_956;
sumr_957<= mulr_1_957 xor mulr_2_957 xor mulr_3_957 xor mulr_4_957;
sumr_958<= mulr_1_958 xor mulr_2_958 xor mulr_3_958 xor mulr_4_958;
sumr_959<= mulr_1_959 xor mulr_2_959 xor mulr_3_959 xor mulr_4_959;
sumr_960<= mulr_1_960 xor mulr_2_960 xor mulr_3_960 xor mulr_4_960;
sumr_961<= mulr_1_961 xor mulr_2_961 xor mulr_3_961 xor mulr_4_961;
sumr_962<= mulr_1_962 xor mulr_2_962 xor mulr_3_962 xor mulr_4_962;
sumr_963<= mulr_1_963 xor mulr_2_963 xor mulr_3_963 xor mulr_4_963;
sumr_964<= mulr_1_964 xor mulr_2_964 xor mulr_3_964 xor mulr_4_964;
sumr_965<= mulr_1_965 xor mulr_2_965 xor mulr_3_965 xor mulr_4_965;
sumr_966<= mulr_1_966 xor mulr_2_966 xor mulr_3_966 xor mulr_4_966;
sumr_967<= mulr_1_967 xor mulr_2_967 xor mulr_3_967 xor mulr_4_967;
sumr_968<= mulr_1_968 xor mulr_2_968 xor mulr_3_968 xor mulr_4_968;
sumr_969<= mulr_1_969 xor mulr_2_969 xor mulr_3_969 xor mulr_4_969;
sumr_970<= mulr_1_970 xor mulr_2_970 xor mulr_3_970 xor mulr_4_970;
sumr_971<= mulr_1_971 xor mulr_2_971 xor mulr_3_971 xor mulr_4_971;
sumr_972<= mulr_1_972 xor mulr_2_972 xor mulr_3_972 xor mulr_4_972;
sumr_973<= mulr_1_973 xor mulr_2_973 xor mulr_3_973 xor mulr_4_973;
sumr_974<= mulr_1_974 xor mulr_2_974 xor mulr_3_974 xor mulr_4_974;
sumr_975<= mulr_1_975 xor mulr_2_975 xor mulr_3_975 xor mulr_4_975;
sumr_976<= mulr_1_976 xor mulr_2_976 xor mulr_3_976 xor mulr_4_976;
sumr_977<= mulr_1_977 xor mulr_2_977 xor mulr_3_977 xor mulr_4_977;
sumr_978<= mulr_1_978 xor mulr_2_978 xor mulr_3_978 xor mulr_4_978;
sumr_979<= mulr_1_979 xor mulr_2_979 xor mulr_3_979 xor mulr_4_979;
sumr_980<= mulr_1_980 xor mulr_2_980 xor mulr_3_980 xor mulr_4_980;
sumr_981<= mulr_1_981 xor mulr_2_981 xor mulr_3_981 xor mulr_4_981;
sumr_982<= mulr_1_982 xor mulr_2_982 xor mulr_3_982 xor mulr_4_982;
sumr_983<= mulr_1_983 xor mulr_2_983 xor mulr_3_983 xor mulr_4_983;
sumr_984<= mulr_1_984 xor mulr_2_984 xor mulr_3_984 xor mulr_4_984;
sumr_985<= mulr_1_985 xor mulr_2_985 xor mulr_3_985 xor mulr_4_985;
sumr_986<= mulr_1_986 xor mulr_2_986 xor mulr_3_986 xor mulr_4_986;
sumr_987<= mulr_1_987 xor mulr_2_987 xor mulr_3_987 xor mulr_4_987;
sumr_988<= mulr_1_988 xor mulr_2_988 xor mulr_3_988 xor mulr_4_988;
sumr_989<= mulr_1_989 xor mulr_2_989 xor mulr_3_989 xor mulr_4_989;
sumr_990<= mulr_1_990 xor mulr_2_990 xor mulr_3_990 xor mulr_4_990;
sumr_991<= mulr_1_991 xor mulr_2_991 xor mulr_3_991 xor mulr_4_991;
sumr_992<= mulr_1_992 xor mulr_2_992 xor mulr_3_992 xor mulr_4_992;
sumr_993<= mulr_1_993 xor mulr_2_993 xor mulr_3_993 xor mulr_4_993;
sumr_994<= mulr_1_994 xor mulr_2_994 xor mulr_3_994 xor mulr_4_994;
sumr_995<= mulr_1_995 xor mulr_2_995 xor mulr_3_995 xor mulr_4_995;
sumr_996<= mulr_1_996 xor mulr_2_996 xor mulr_3_996 xor mulr_4_996;
sumr_997<= mulr_1_997 xor mulr_2_997 xor mulr_3_997 xor mulr_4_997;
sumr_998<= mulr_1_998 xor mulr_2_998 xor mulr_3_998 xor mulr_4_998;
sumr_999<= mulr_1_999 xor mulr_2_999 xor mulr_3_999 xor mulr_4_999;
sumr_1000<= mulr_1_1000 xor mulr_2_1000 xor mulr_3_1000 xor mulr_4_1000;
sumr_1001<= mulr_1_1001 xor mulr_2_1001 xor mulr_3_1001 xor mulr_4_1001;
sumr_1002<= mulr_1_1002 xor mulr_2_1002 xor mulr_3_1002 xor mulr_4_1002;
sumr_1003<= mulr_1_1003 xor mulr_2_1003 xor mulr_3_1003 xor mulr_4_1003;
sumr_1004<= mulr_1_1004 xor mulr_2_1004 xor mulr_3_1004 xor mulr_4_1004;
sumr_1005<= mulr_1_1005 xor mulr_2_1005 xor mulr_3_1005 xor mulr_4_1005;
sumr_1006<= mulr_1_1006 xor mulr_2_1006 xor mulr_3_1006 xor mulr_4_1006;
sumr_1007<= mulr_1_1007 xor mulr_2_1007 xor mulr_3_1007 xor mulr_4_1007;
sumr_1008<= mulr_1_1008 xor mulr_2_1008 xor mulr_3_1008 xor mulr_4_1008;
sumr_1009<= mulr_1_1009 xor mulr_2_1009 xor mulr_3_1009 xor mulr_4_1009;
sumr_1010<= mulr_1_1010 xor mulr_2_1010 xor mulr_3_1010 xor mulr_4_1010;
sumr_1011<= mulr_1_1011 xor mulr_2_1011 xor mulr_3_1011 xor mulr_4_1011;
sumr_1012<= mulr_1_1012 xor mulr_2_1012 xor mulr_3_1012 xor mulr_4_1012;
sumr_1013<= mulr_1_1013 xor mulr_2_1013 xor mulr_3_1013 xor mulr_4_1013;
sumr_1014<= mulr_1_1014 xor mulr_2_1014 xor mulr_3_1014 xor mulr_4_1014;
sumr_1015<= mulr_1_1015 xor mulr_2_1015 xor mulr_3_1015 xor mulr_4_1015;
sumr_1016<= mulr_1_1016 xor mulr_2_1016 xor mulr_3_1016 xor mulr_4_1016;
sumr_1017<= mulr_1_1017 xor mulr_2_1017 xor mulr_3_1017 xor mulr_4_1017;
sumr_1018<= mulr_1_1018 xor mulr_2_1018 xor mulr_3_1018 xor mulr_4_1018;
sumr_1019<= mulr_1_1019 xor mulr_2_1019 xor mulr_3_1019 xor mulr_4_1019;
sumr_1020<= mulr_1_1020 xor mulr_2_1020 xor mulr_3_1020 xor mulr_4_1020;
sumr_1021<= mulr_1_1021 xor mulr_2_1021 xor mulr_3_1021 xor mulr_4_1021;
sumr_1022<= mulr_1_1022 xor mulr_2_1022 xor mulr_3_1022 xor mulr_4_1022;
sumr_1023<= mulr_1_1023 xor mulr_2_1023 xor mulr_3_1023 xor mulr_4_1023;
E(1022)<=not ( sumr_1(0) or sumr_1(1) or sumr_1(2) or sumr_1(3) or sumr_1(4) or sumr_1(5) or sumr_1(6) or sumr_1(7) or sumr_1(8) or sumr_1(9));
E(1021)<=not ( sumr_2(0) or sumr_2(1) or sumr_2(2) or sumr_2(3) or sumr_2(4) or sumr_2(5) or sumr_2(6) or sumr_2(7) or sumr_2(8) or sumr_2(9));
E(1020)<=not ( sumr_3(0) or sumr_3(1) or sumr_3(2) or sumr_3(3) or sumr_3(4) or sumr_3(5) or sumr_3(6) or sumr_3(7) or sumr_3(8) or sumr_3(9));
E(1019)<=not ( sumr_4(0) or sumr_4(1) or sumr_4(2) or sumr_4(3) or sumr_4(4) or sumr_4(5) or sumr_4(6) or sumr_4(7) or sumr_4(8) or sumr_4(9));
E(1018)<=not ( sumr_5(0) or sumr_5(1) or sumr_5(2) or sumr_5(3) or sumr_5(4) or sumr_5(5) or sumr_5(6) or sumr_5(7) or sumr_5(8) or sumr_5(9));
E(1017)<=not ( sumr_6(0) or sumr_6(1) or sumr_6(2) or sumr_6(3) or sumr_6(4) or sumr_6(5) or sumr_6(6) or sumr_6(7) or sumr_6(8) or sumr_6(9));
E(1016)<=not ( sumr_7(0) or sumr_7(1) or sumr_7(2) or sumr_7(3) or sumr_7(4) or sumr_7(5) or sumr_7(6) or sumr_7(7) or sumr_7(8) or sumr_7(9));
E(1015)<=not ( sumr_8(0) or sumr_8(1) or sumr_8(2) or sumr_8(3) or sumr_8(4) or sumr_8(5) or sumr_8(6) or sumr_8(7) or sumr_8(8) or sumr_8(9));
E(1014)<=not ( sumr_9(0) or sumr_9(1) or sumr_9(2) or sumr_9(3) or sumr_9(4) or sumr_9(5) or sumr_9(6) or sumr_9(7) or sumr_9(8) or sumr_9(9));
E(1013)<=not ( sumr_10(0) or sumr_10(1) or sumr_10(2) or sumr_10(3) or sumr_10(4) or sumr_10(5) or sumr_10(6) or sumr_10(7) or sumr_10(8) or sumr_10(9));
E(1012)<=not ( sumr_11(0) or sumr_11(1) or sumr_11(2) or sumr_11(3) or sumr_11(4) or sumr_11(5) or sumr_11(6) or sumr_11(7) or sumr_11(8) or sumr_11(9));
E(1011)<=not ( sumr_12(0) or sumr_12(1) or sumr_12(2) or sumr_12(3) or sumr_12(4) or sumr_12(5) or sumr_12(6) or sumr_12(7) or sumr_12(8) or sumr_12(9));
E(1010)<=not ( sumr_13(0) or sumr_13(1) or sumr_13(2) or sumr_13(3) or sumr_13(4) or sumr_13(5) or sumr_13(6) or sumr_13(7) or sumr_13(8) or sumr_13(9));
E(1009)<=not ( sumr_14(0) or sumr_14(1) or sumr_14(2) or sumr_14(3) or sumr_14(4) or sumr_14(5) or sumr_14(6) or sumr_14(7) or sumr_14(8) or sumr_14(9));
E(1008)<=not ( sumr_15(0) or sumr_15(1) or sumr_15(2) or sumr_15(3) or sumr_15(4) or sumr_15(5) or sumr_15(6) or sumr_15(7) or sumr_15(8) or sumr_15(9));
E(1007)<=not ( sumr_16(0) or sumr_16(1) or sumr_16(2) or sumr_16(3) or sumr_16(4) or sumr_16(5) or sumr_16(6) or sumr_16(7) or sumr_16(8) or sumr_16(9));
E(1006)<=not ( sumr_17(0) or sumr_17(1) or sumr_17(2) or sumr_17(3) or sumr_17(4) or sumr_17(5) or sumr_17(6) or sumr_17(7) or sumr_17(8) or sumr_17(9));
E(1005)<=not ( sumr_18(0) or sumr_18(1) or sumr_18(2) or sumr_18(3) or sumr_18(4) or sumr_18(5) or sumr_18(6) or sumr_18(7) or sumr_18(8) or sumr_18(9));
E(1004)<=not ( sumr_19(0) or sumr_19(1) or sumr_19(2) or sumr_19(3) or sumr_19(4) or sumr_19(5) or sumr_19(6) or sumr_19(7) or sumr_19(8) or sumr_19(9));
E(1003)<=not ( sumr_20(0) or sumr_20(1) or sumr_20(2) or sumr_20(3) or sumr_20(4) or sumr_20(5) or sumr_20(6) or sumr_20(7) or sumr_20(8) or sumr_20(9));
E(1002)<=not ( sumr_21(0) or sumr_21(1) or sumr_21(2) or sumr_21(3) or sumr_21(4) or sumr_21(5) or sumr_21(6) or sumr_21(7) or sumr_21(8) or sumr_21(9));
E(1001)<=not ( sumr_22(0) or sumr_22(1) or sumr_22(2) or sumr_22(3) or sumr_22(4) or sumr_22(5) or sumr_22(6) or sumr_22(7) or sumr_22(8) or sumr_22(9));
E(1000)<=not ( sumr_23(0) or sumr_23(1) or sumr_23(2) or sumr_23(3) or sumr_23(4) or sumr_23(5) or sumr_23(6) or sumr_23(7) or sumr_23(8) or sumr_23(9));
E(999)<=not ( sumr_24(0) or sumr_24(1) or sumr_24(2) or sumr_24(3) or sumr_24(4) or sumr_24(5) or sumr_24(6) or sumr_24(7) or sumr_24(8) or sumr_24(9));
E(998)<=not ( sumr_25(0) or sumr_25(1) or sumr_25(2) or sumr_25(3) or sumr_25(4) or sumr_25(5) or sumr_25(6) or sumr_25(7) or sumr_25(8) or sumr_25(9));
E(997)<=not ( sumr_26(0) or sumr_26(1) or sumr_26(2) or sumr_26(3) or sumr_26(4) or sumr_26(5) or sumr_26(6) or sumr_26(7) or sumr_26(8) or sumr_26(9));
E(996)<=not ( sumr_27(0) or sumr_27(1) or sumr_27(2) or sumr_27(3) or sumr_27(4) or sumr_27(5) or sumr_27(6) or sumr_27(7) or sumr_27(8) or sumr_27(9));
E(995)<=not ( sumr_28(0) or sumr_28(1) or sumr_28(2) or sumr_28(3) or sumr_28(4) or sumr_28(5) or sumr_28(6) or sumr_28(7) or sumr_28(8) or sumr_28(9));
E(994)<=not ( sumr_29(0) or sumr_29(1) or sumr_29(2) or sumr_29(3) or sumr_29(4) or sumr_29(5) or sumr_29(6) or sumr_29(7) or sumr_29(8) or sumr_29(9));
E(993)<=not ( sumr_30(0) or sumr_30(1) or sumr_30(2) or sumr_30(3) or sumr_30(4) or sumr_30(5) or sumr_30(6) or sumr_30(7) or sumr_30(8) or sumr_30(9));
E(992)<=not ( sumr_31(0) or sumr_31(1) or sumr_31(2) or sumr_31(3) or sumr_31(4) or sumr_31(5) or sumr_31(6) or sumr_31(7) or sumr_31(8) or sumr_31(9));
E(991)<=not ( sumr_32(0) or sumr_32(1) or sumr_32(2) or sumr_32(3) or sumr_32(4) or sumr_32(5) or sumr_32(6) or sumr_32(7) or sumr_32(8) or sumr_32(9));
E(990)<=not ( sumr_33(0) or sumr_33(1) or sumr_33(2) or sumr_33(3) or sumr_33(4) or sumr_33(5) or sumr_33(6) or sumr_33(7) or sumr_33(8) or sumr_33(9));
E(989)<=not ( sumr_34(0) or sumr_34(1) or sumr_34(2) or sumr_34(3) or sumr_34(4) or sumr_34(5) or sumr_34(6) or sumr_34(7) or sumr_34(8) or sumr_34(9));
E(988)<=not ( sumr_35(0) or sumr_35(1) or sumr_35(2) or sumr_35(3) or sumr_35(4) or sumr_35(5) or sumr_35(6) or sumr_35(7) or sumr_35(8) or sumr_35(9));
E(987)<=not ( sumr_36(0) or sumr_36(1) or sumr_36(2) or sumr_36(3) or sumr_36(4) or sumr_36(5) or sumr_36(6) or sumr_36(7) or sumr_36(8) or sumr_36(9));
E(986)<=not ( sumr_37(0) or sumr_37(1) or sumr_37(2) or sumr_37(3) or sumr_37(4) or sumr_37(5) or sumr_37(6) or sumr_37(7) or sumr_37(8) or sumr_37(9));
E(985)<=not ( sumr_38(0) or sumr_38(1) or sumr_38(2) or sumr_38(3) or sumr_38(4) or sumr_38(5) or sumr_38(6) or sumr_38(7) or sumr_38(8) or sumr_38(9));
E(984)<=not ( sumr_39(0) or sumr_39(1) or sumr_39(2) or sumr_39(3) or sumr_39(4) or sumr_39(5) or sumr_39(6) or sumr_39(7) or sumr_39(8) or sumr_39(9));
E(983)<=not ( sumr_40(0) or sumr_40(1) or sumr_40(2) or sumr_40(3) or sumr_40(4) or sumr_40(5) or sumr_40(6) or sumr_40(7) or sumr_40(8) or sumr_40(9));
E(982)<=not ( sumr_41(0) or sumr_41(1) or sumr_41(2) or sumr_41(3) or sumr_41(4) or sumr_41(5) or sumr_41(6) or sumr_41(7) or sumr_41(8) or sumr_41(9));
E(981)<=not ( sumr_42(0) or sumr_42(1) or sumr_42(2) or sumr_42(3) or sumr_42(4) or sumr_42(5) or sumr_42(6) or sumr_42(7) or sumr_42(8) or sumr_42(9));
E(980)<=not ( sumr_43(0) or sumr_43(1) or sumr_43(2) or sumr_43(3) or sumr_43(4) or sumr_43(5) or sumr_43(6) or sumr_43(7) or sumr_43(8) or sumr_43(9));
E(979)<=not ( sumr_44(0) or sumr_44(1) or sumr_44(2) or sumr_44(3) or sumr_44(4) or sumr_44(5) or sumr_44(6) or sumr_44(7) or sumr_44(8) or sumr_44(9));
E(978)<=not ( sumr_45(0) or sumr_45(1) or sumr_45(2) or sumr_45(3) or sumr_45(4) or sumr_45(5) or sumr_45(6) or sumr_45(7) or sumr_45(8) or sumr_45(9));
E(977)<=not ( sumr_46(0) or sumr_46(1) or sumr_46(2) or sumr_46(3) or sumr_46(4) or sumr_46(5) or sumr_46(6) or sumr_46(7) or sumr_46(8) or sumr_46(9));
E(976)<=not ( sumr_47(0) or sumr_47(1) or sumr_47(2) or sumr_47(3) or sumr_47(4) or sumr_47(5) or sumr_47(6) or sumr_47(7) or sumr_47(8) or sumr_47(9));
E(975)<=not ( sumr_48(0) or sumr_48(1) or sumr_48(2) or sumr_48(3) or sumr_48(4) or sumr_48(5) or sumr_48(6) or sumr_48(7) or sumr_48(8) or sumr_48(9));
E(974)<=not ( sumr_49(0) or sumr_49(1) or sumr_49(2) or sumr_49(3) or sumr_49(4) or sumr_49(5) or sumr_49(6) or sumr_49(7) or sumr_49(8) or sumr_49(9));
E(973)<=not ( sumr_50(0) or sumr_50(1) or sumr_50(2) or sumr_50(3) or sumr_50(4) or sumr_50(5) or sumr_50(6) or sumr_50(7) or sumr_50(8) or sumr_50(9));
E(972)<=not ( sumr_51(0) or sumr_51(1) or sumr_51(2) or sumr_51(3) or sumr_51(4) or sumr_51(5) or sumr_51(6) or sumr_51(7) or sumr_51(8) or sumr_51(9));
E(971)<=not ( sumr_52(0) or sumr_52(1) or sumr_52(2) or sumr_52(3) or sumr_52(4) or sumr_52(5) or sumr_52(6) or sumr_52(7) or sumr_52(8) or sumr_52(9));
E(970)<=not ( sumr_53(0) or sumr_53(1) or sumr_53(2) or sumr_53(3) or sumr_53(4) or sumr_53(5) or sumr_53(6) or sumr_53(7) or sumr_53(8) or sumr_53(9));
E(969)<=not ( sumr_54(0) or sumr_54(1) or sumr_54(2) or sumr_54(3) or sumr_54(4) or sumr_54(5) or sumr_54(6) or sumr_54(7) or sumr_54(8) or sumr_54(9));
E(968)<=not ( sumr_55(0) or sumr_55(1) or sumr_55(2) or sumr_55(3) or sumr_55(4) or sumr_55(5) or sumr_55(6) or sumr_55(7) or sumr_55(8) or sumr_55(9));
E(967)<=not ( sumr_56(0) or sumr_56(1) or sumr_56(2) or sumr_56(3) or sumr_56(4) or sumr_56(5) or sumr_56(6) or sumr_56(7) or sumr_56(8) or sumr_56(9));
E(966)<=not ( sumr_57(0) or sumr_57(1) or sumr_57(2) or sumr_57(3) or sumr_57(4) or sumr_57(5) or sumr_57(6) or sumr_57(7) or sumr_57(8) or sumr_57(9));
E(965)<=not ( sumr_58(0) or sumr_58(1) or sumr_58(2) or sumr_58(3) or sumr_58(4) or sumr_58(5) or sumr_58(6) or sumr_58(7) or sumr_58(8) or sumr_58(9));
E(964)<=not ( sumr_59(0) or sumr_59(1) or sumr_59(2) or sumr_59(3) or sumr_59(4) or sumr_59(5) or sumr_59(6) or sumr_59(7) or sumr_59(8) or sumr_59(9));
E(963)<=not ( sumr_60(0) or sumr_60(1) or sumr_60(2) or sumr_60(3) or sumr_60(4) or sumr_60(5) or sumr_60(6) or sumr_60(7) or sumr_60(8) or sumr_60(9));
E(962)<=not ( sumr_61(0) or sumr_61(1) or sumr_61(2) or sumr_61(3) or sumr_61(4) or sumr_61(5) or sumr_61(6) or sumr_61(7) or sumr_61(8) or sumr_61(9));
E(961)<=not ( sumr_62(0) or sumr_62(1) or sumr_62(2) or sumr_62(3) or sumr_62(4) or sumr_62(5) or sumr_62(6) or sumr_62(7) or sumr_62(8) or sumr_62(9));
E(960)<=not ( sumr_63(0) or sumr_63(1) or sumr_63(2) or sumr_63(3) or sumr_63(4) or sumr_63(5) or sumr_63(6) or sumr_63(7) or sumr_63(8) or sumr_63(9));
E(959)<=not ( sumr_64(0) or sumr_64(1) or sumr_64(2) or sumr_64(3) or sumr_64(4) or sumr_64(5) or sumr_64(6) or sumr_64(7) or sumr_64(8) or sumr_64(9));
E(958)<=not ( sumr_65(0) or sumr_65(1) or sumr_65(2) or sumr_65(3) or sumr_65(4) or sumr_65(5) or sumr_65(6) or sumr_65(7) or sumr_65(8) or sumr_65(9));
E(957)<=not ( sumr_66(0) or sumr_66(1) or sumr_66(2) or sumr_66(3) or sumr_66(4) or sumr_66(5) or sumr_66(6) or sumr_66(7) or sumr_66(8) or sumr_66(9));
E(956)<=not ( sumr_67(0) or sumr_67(1) or sumr_67(2) or sumr_67(3) or sumr_67(4) or sumr_67(5) or sumr_67(6) or sumr_67(7) or sumr_67(8) or sumr_67(9));
E(955)<=not ( sumr_68(0) or sumr_68(1) or sumr_68(2) or sumr_68(3) or sumr_68(4) or sumr_68(5) or sumr_68(6) or sumr_68(7) or sumr_68(8) or sumr_68(9));
E(954)<=not ( sumr_69(0) or sumr_69(1) or sumr_69(2) or sumr_69(3) or sumr_69(4) or sumr_69(5) or sumr_69(6) or sumr_69(7) or sumr_69(8) or sumr_69(9));
E(953)<=not ( sumr_70(0) or sumr_70(1) or sumr_70(2) or sumr_70(3) or sumr_70(4) or sumr_70(5) or sumr_70(6) or sumr_70(7) or sumr_70(8) or sumr_70(9));
E(952)<=not ( sumr_71(0) or sumr_71(1) or sumr_71(2) or sumr_71(3) or sumr_71(4) or sumr_71(5) or sumr_71(6) or sumr_71(7) or sumr_71(8) or sumr_71(9));
E(951)<=not ( sumr_72(0) or sumr_72(1) or sumr_72(2) or sumr_72(3) or sumr_72(4) or sumr_72(5) or sumr_72(6) or sumr_72(7) or sumr_72(8) or sumr_72(9));
E(950)<=not ( sumr_73(0) or sumr_73(1) or sumr_73(2) or sumr_73(3) or sumr_73(4) or sumr_73(5) or sumr_73(6) or sumr_73(7) or sumr_73(8) or sumr_73(9));
E(949)<=not ( sumr_74(0) or sumr_74(1) or sumr_74(2) or sumr_74(3) or sumr_74(4) or sumr_74(5) or sumr_74(6) or sumr_74(7) or sumr_74(8) or sumr_74(9));
E(948)<=not ( sumr_75(0) or sumr_75(1) or sumr_75(2) or sumr_75(3) or sumr_75(4) or sumr_75(5) or sumr_75(6) or sumr_75(7) or sumr_75(8) or sumr_75(9));
E(947)<=not ( sumr_76(0) or sumr_76(1) or sumr_76(2) or sumr_76(3) or sumr_76(4) or sumr_76(5) or sumr_76(6) or sumr_76(7) or sumr_76(8) or sumr_76(9));
E(946)<=not ( sumr_77(0) or sumr_77(1) or sumr_77(2) or sumr_77(3) or sumr_77(4) or sumr_77(5) or sumr_77(6) or sumr_77(7) or sumr_77(8) or sumr_77(9));
E(945)<=not ( sumr_78(0) or sumr_78(1) or sumr_78(2) or sumr_78(3) or sumr_78(4) or sumr_78(5) or sumr_78(6) or sumr_78(7) or sumr_78(8) or sumr_78(9));
E(944)<=not ( sumr_79(0) or sumr_79(1) or sumr_79(2) or sumr_79(3) or sumr_79(4) or sumr_79(5) or sumr_79(6) or sumr_79(7) or sumr_79(8) or sumr_79(9));
E(943)<=not ( sumr_80(0) or sumr_80(1) or sumr_80(2) or sumr_80(3) or sumr_80(4) or sumr_80(5) or sumr_80(6) or sumr_80(7) or sumr_80(8) or sumr_80(9));
E(942)<=not ( sumr_81(0) or sumr_81(1) or sumr_81(2) or sumr_81(3) or sumr_81(4) or sumr_81(5) or sumr_81(6) or sumr_81(7) or sumr_81(8) or sumr_81(9));
E(941)<=not ( sumr_82(0) or sumr_82(1) or sumr_82(2) or sumr_82(3) or sumr_82(4) or sumr_82(5) or sumr_82(6) or sumr_82(7) or sumr_82(8) or sumr_82(9));
E(940)<=not ( sumr_83(0) or sumr_83(1) or sumr_83(2) or sumr_83(3) or sumr_83(4) or sumr_83(5) or sumr_83(6) or sumr_83(7) or sumr_83(8) or sumr_83(9));
E(939)<=not ( sumr_84(0) or sumr_84(1) or sumr_84(2) or sumr_84(3) or sumr_84(4) or sumr_84(5) or sumr_84(6) or sumr_84(7) or sumr_84(8) or sumr_84(9));
E(938)<=not ( sumr_85(0) or sumr_85(1) or sumr_85(2) or sumr_85(3) or sumr_85(4) or sumr_85(5) or sumr_85(6) or sumr_85(7) or sumr_85(8) or sumr_85(9));
E(937)<=not ( sumr_86(0) or sumr_86(1) or sumr_86(2) or sumr_86(3) or sumr_86(4) or sumr_86(5) or sumr_86(6) or sumr_86(7) or sumr_86(8) or sumr_86(9));
E(936)<=not ( sumr_87(0) or sumr_87(1) or sumr_87(2) or sumr_87(3) or sumr_87(4) or sumr_87(5) or sumr_87(6) or sumr_87(7) or sumr_87(8) or sumr_87(9));
E(935)<=not ( sumr_88(0) or sumr_88(1) or sumr_88(2) or sumr_88(3) or sumr_88(4) or sumr_88(5) or sumr_88(6) or sumr_88(7) or sumr_88(8) or sumr_88(9));
E(934)<=not ( sumr_89(0) or sumr_89(1) or sumr_89(2) or sumr_89(3) or sumr_89(4) or sumr_89(5) or sumr_89(6) or sumr_89(7) or sumr_89(8) or sumr_89(9));
E(933)<=not ( sumr_90(0) or sumr_90(1) or sumr_90(2) or sumr_90(3) or sumr_90(4) or sumr_90(5) or sumr_90(6) or sumr_90(7) or sumr_90(8) or sumr_90(9));
E(932)<=not ( sumr_91(0) or sumr_91(1) or sumr_91(2) or sumr_91(3) or sumr_91(4) or sumr_91(5) or sumr_91(6) or sumr_91(7) or sumr_91(8) or sumr_91(9));
E(931)<=not ( sumr_92(0) or sumr_92(1) or sumr_92(2) or sumr_92(3) or sumr_92(4) or sumr_92(5) or sumr_92(6) or sumr_92(7) or sumr_92(8) or sumr_92(9));
E(930)<=not ( sumr_93(0) or sumr_93(1) or sumr_93(2) or sumr_93(3) or sumr_93(4) or sumr_93(5) or sumr_93(6) or sumr_93(7) or sumr_93(8) or sumr_93(9));
E(929)<=not ( sumr_94(0) or sumr_94(1) or sumr_94(2) or sumr_94(3) or sumr_94(4) or sumr_94(5) or sumr_94(6) or sumr_94(7) or sumr_94(8) or sumr_94(9));
E(928)<=not ( sumr_95(0) or sumr_95(1) or sumr_95(2) or sumr_95(3) or sumr_95(4) or sumr_95(5) or sumr_95(6) or sumr_95(7) or sumr_95(8) or sumr_95(9));
E(927)<=not ( sumr_96(0) or sumr_96(1) or sumr_96(2) or sumr_96(3) or sumr_96(4) or sumr_96(5) or sumr_96(6) or sumr_96(7) or sumr_96(8) or sumr_96(9));
E(926)<=not ( sumr_97(0) or sumr_97(1) or sumr_97(2) or sumr_97(3) or sumr_97(4) or sumr_97(5) or sumr_97(6) or sumr_97(7) or sumr_97(8) or sumr_97(9));
E(925)<=not ( sumr_98(0) or sumr_98(1) or sumr_98(2) or sumr_98(3) or sumr_98(4) or sumr_98(5) or sumr_98(6) or sumr_98(7) or sumr_98(8) or sumr_98(9));
E(924)<=not ( sumr_99(0) or sumr_99(1) or sumr_99(2) or sumr_99(3) or sumr_99(4) or sumr_99(5) or sumr_99(6) or sumr_99(7) or sumr_99(8) or sumr_99(9));
E(923)<=not ( sumr_100(0) or sumr_100(1) or sumr_100(2) or sumr_100(3) or sumr_100(4) or sumr_100(5) or sumr_100(6) or sumr_100(7) or sumr_100(8) or sumr_100(9));
E(922)<=not ( sumr_101(0) or sumr_101(1) or sumr_101(2) or sumr_101(3) or sumr_101(4) or sumr_101(5) or sumr_101(6) or sumr_101(7) or sumr_101(8) or sumr_101(9));
E(921)<=not ( sumr_102(0) or sumr_102(1) or sumr_102(2) or sumr_102(3) or sumr_102(4) or sumr_102(5) or sumr_102(6) or sumr_102(7) or sumr_102(8) or sumr_102(9));
E(920)<=not ( sumr_103(0) or sumr_103(1) or sumr_103(2) or sumr_103(3) or sumr_103(4) or sumr_103(5) or sumr_103(6) or sumr_103(7) or sumr_103(8) or sumr_103(9));
E(919)<=not ( sumr_104(0) or sumr_104(1) or sumr_104(2) or sumr_104(3) or sumr_104(4) or sumr_104(5) or sumr_104(6) or sumr_104(7) or sumr_104(8) or sumr_104(9));
E(918)<=not ( sumr_105(0) or sumr_105(1) or sumr_105(2) or sumr_105(3) or sumr_105(4) or sumr_105(5) or sumr_105(6) or sumr_105(7) or sumr_105(8) or sumr_105(9));
E(917)<=not ( sumr_106(0) or sumr_106(1) or sumr_106(2) or sumr_106(3) or sumr_106(4) or sumr_106(5) or sumr_106(6) or sumr_106(7) or sumr_106(8) or sumr_106(9));
E(916)<=not ( sumr_107(0) or sumr_107(1) or sumr_107(2) or sumr_107(3) or sumr_107(4) or sumr_107(5) or sumr_107(6) or sumr_107(7) or sumr_107(8) or sumr_107(9));
E(915)<=not ( sumr_108(0) or sumr_108(1) or sumr_108(2) or sumr_108(3) or sumr_108(4) or sumr_108(5) or sumr_108(6) or sumr_108(7) or sumr_108(8) or sumr_108(9));
E(914)<=not ( sumr_109(0) or sumr_109(1) or sumr_109(2) or sumr_109(3) or sumr_109(4) or sumr_109(5) or sumr_109(6) or sumr_109(7) or sumr_109(8) or sumr_109(9));
E(913)<=not ( sumr_110(0) or sumr_110(1) or sumr_110(2) or sumr_110(3) or sumr_110(4) or sumr_110(5) or sumr_110(6) or sumr_110(7) or sumr_110(8) or sumr_110(9));
E(912)<=not ( sumr_111(0) or sumr_111(1) or sumr_111(2) or sumr_111(3) or sumr_111(4) or sumr_111(5) or sumr_111(6) or sumr_111(7) or sumr_111(8) or sumr_111(9));
E(911)<=not ( sumr_112(0) or sumr_112(1) or sumr_112(2) or sumr_112(3) or sumr_112(4) or sumr_112(5) or sumr_112(6) or sumr_112(7) or sumr_112(8) or sumr_112(9));
E(910)<=not ( sumr_113(0) or sumr_113(1) or sumr_113(2) or sumr_113(3) or sumr_113(4) or sumr_113(5) or sumr_113(6) or sumr_113(7) or sumr_113(8) or sumr_113(9));
E(909)<=not ( sumr_114(0) or sumr_114(1) or sumr_114(2) or sumr_114(3) or sumr_114(4) or sumr_114(5) or sumr_114(6) or sumr_114(7) or sumr_114(8) or sumr_114(9));
E(908)<=not ( sumr_115(0) or sumr_115(1) or sumr_115(2) or sumr_115(3) or sumr_115(4) or sumr_115(5) or sumr_115(6) or sumr_115(7) or sumr_115(8) or sumr_115(9));
E(907)<=not ( sumr_116(0) or sumr_116(1) or sumr_116(2) or sumr_116(3) or sumr_116(4) or sumr_116(5) or sumr_116(6) or sumr_116(7) or sumr_116(8) or sumr_116(9));
E(906)<=not ( sumr_117(0) or sumr_117(1) or sumr_117(2) or sumr_117(3) or sumr_117(4) or sumr_117(5) or sumr_117(6) or sumr_117(7) or sumr_117(8) or sumr_117(9));
E(905)<=not ( sumr_118(0) or sumr_118(1) or sumr_118(2) or sumr_118(3) or sumr_118(4) or sumr_118(5) or sumr_118(6) or sumr_118(7) or sumr_118(8) or sumr_118(9));
E(904)<=not ( sumr_119(0) or sumr_119(1) or sumr_119(2) or sumr_119(3) or sumr_119(4) or sumr_119(5) or sumr_119(6) or sumr_119(7) or sumr_119(8) or sumr_119(9));
E(903)<=not ( sumr_120(0) or sumr_120(1) or sumr_120(2) or sumr_120(3) or sumr_120(4) or sumr_120(5) or sumr_120(6) or sumr_120(7) or sumr_120(8) or sumr_120(9));
E(902)<=not ( sumr_121(0) or sumr_121(1) or sumr_121(2) or sumr_121(3) or sumr_121(4) or sumr_121(5) or sumr_121(6) or sumr_121(7) or sumr_121(8) or sumr_121(9));
E(901)<=not ( sumr_122(0) or sumr_122(1) or sumr_122(2) or sumr_122(3) or sumr_122(4) or sumr_122(5) or sumr_122(6) or sumr_122(7) or sumr_122(8) or sumr_122(9));
E(900)<=not ( sumr_123(0) or sumr_123(1) or sumr_123(2) or sumr_123(3) or sumr_123(4) or sumr_123(5) or sumr_123(6) or sumr_123(7) or sumr_123(8) or sumr_123(9));
E(899)<=not ( sumr_124(0) or sumr_124(1) or sumr_124(2) or sumr_124(3) or sumr_124(4) or sumr_124(5) or sumr_124(6) or sumr_124(7) or sumr_124(8) or sumr_124(9));
E(898)<=not ( sumr_125(0) or sumr_125(1) or sumr_125(2) or sumr_125(3) or sumr_125(4) or sumr_125(5) or sumr_125(6) or sumr_125(7) or sumr_125(8) or sumr_125(9));
E(897)<=not ( sumr_126(0) or sumr_126(1) or sumr_126(2) or sumr_126(3) or sumr_126(4) or sumr_126(5) or sumr_126(6) or sumr_126(7) or sumr_126(8) or sumr_126(9));
E(896)<=not ( sumr_127(0) or sumr_127(1) or sumr_127(2) or sumr_127(3) or sumr_127(4) or sumr_127(5) or sumr_127(6) or sumr_127(7) or sumr_127(8) or sumr_127(9));
E(895)<=not ( sumr_128(0) or sumr_128(1) or sumr_128(2) or sumr_128(3) or sumr_128(4) or sumr_128(5) or sumr_128(6) or sumr_128(7) or sumr_128(8) or sumr_128(9));
E(894)<=not ( sumr_129(0) or sumr_129(1) or sumr_129(2) or sumr_129(3) or sumr_129(4) or sumr_129(5) or sumr_129(6) or sumr_129(7) or sumr_129(8) or sumr_129(9));
E(893)<=not ( sumr_130(0) or sumr_130(1) or sumr_130(2) or sumr_130(3) or sumr_130(4) or sumr_130(5) or sumr_130(6) or sumr_130(7) or sumr_130(8) or sumr_130(9));
E(892)<=not ( sumr_131(0) or sumr_131(1) or sumr_131(2) or sumr_131(3) or sumr_131(4) or sumr_131(5) or sumr_131(6) or sumr_131(7) or sumr_131(8) or sumr_131(9));
E(891)<=not ( sumr_132(0) or sumr_132(1) or sumr_132(2) or sumr_132(3) or sumr_132(4) or sumr_132(5) or sumr_132(6) or sumr_132(7) or sumr_132(8) or sumr_132(9));
E(890)<=not ( sumr_133(0) or sumr_133(1) or sumr_133(2) or sumr_133(3) or sumr_133(4) or sumr_133(5) or sumr_133(6) or sumr_133(7) or sumr_133(8) or sumr_133(9));
E(889)<=not ( sumr_134(0) or sumr_134(1) or sumr_134(2) or sumr_134(3) or sumr_134(4) or sumr_134(5) or sumr_134(6) or sumr_134(7) or sumr_134(8) or sumr_134(9));
E(888)<=not ( sumr_135(0) or sumr_135(1) or sumr_135(2) or sumr_135(3) or sumr_135(4) or sumr_135(5) or sumr_135(6) or sumr_135(7) or sumr_135(8) or sumr_135(9));
E(887)<=not ( sumr_136(0) or sumr_136(1) or sumr_136(2) or sumr_136(3) or sumr_136(4) or sumr_136(5) or sumr_136(6) or sumr_136(7) or sumr_136(8) or sumr_136(9));
E(886)<=not ( sumr_137(0) or sumr_137(1) or sumr_137(2) or sumr_137(3) or sumr_137(4) or sumr_137(5) or sumr_137(6) or sumr_137(7) or sumr_137(8) or sumr_137(9));
E(885)<=not ( sumr_138(0) or sumr_138(1) or sumr_138(2) or sumr_138(3) or sumr_138(4) or sumr_138(5) or sumr_138(6) or sumr_138(7) or sumr_138(8) or sumr_138(9));
E(884)<=not ( sumr_139(0) or sumr_139(1) or sumr_139(2) or sumr_139(3) or sumr_139(4) or sumr_139(5) or sumr_139(6) or sumr_139(7) or sumr_139(8) or sumr_139(9));
E(883)<=not ( sumr_140(0) or sumr_140(1) or sumr_140(2) or sumr_140(3) or sumr_140(4) or sumr_140(5) or sumr_140(6) or sumr_140(7) or sumr_140(8) or sumr_140(9));
E(882)<=not ( sumr_141(0) or sumr_141(1) or sumr_141(2) or sumr_141(3) or sumr_141(4) or sumr_141(5) or sumr_141(6) or sumr_141(7) or sumr_141(8) or sumr_141(9));
E(881)<=not ( sumr_142(0) or sumr_142(1) or sumr_142(2) or sumr_142(3) or sumr_142(4) or sumr_142(5) or sumr_142(6) or sumr_142(7) or sumr_142(8) or sumr_142(9));
E(880)<=not ( sumr_143(0) or sumr_143(1) or sumr_143(2) or sumr_143(3) or sumr_143(4) or sumr_143(5) or sumr_143(6) or sumr_143(7) or sumr_143(8) or sumr_143(9));
E(879)<=not ( sumr_144(0) or sumr_144(1) or sumr_144(2) or sumr_144(3) or sumr_144(4) or sumr_144(5) or sumr_144(6) or sumr_144(7) or sumr_144(8) or sumr_144(9));
E(878)<=not ( sumr_145(0) or sumr_145(1) or sumr_145(2) or sumr_145(3) or sumr_145(4) or sumr_145(5) or sumr_145(6) or sumr_145(7) or sumr_145(8) or sumr_145(9));
E(877)<=not ( sumr_146(0) or sumr_146(1) or sumr_146(2) or sumr_146(3) or sumr_146(4) or sumr_146(5) or sumr_146(6) or sumr_146(7) or sumr_146(8) or sumr_146(9));
E(876)<=not ( sumr_147(0) or sumr_147(1) or sumr_147(2) or sumr_147(3) or sumr_147(4) or sumr_147(5) or sumr_147(6) or sumr_147(7) or sumr_147(8) or sumr_147(9));
E(875)<=not ( sumr_148(0) or sumr_148(1) or sumr_148(2) or sumr_148(3) or sumr_148(4) or sumr_148(5) or sumr_148(6) or sumr_148(7) or sumr_148(8) or sumr_148(9));
E(874)<=not ( sumr_149(0) or sumr_149(1) or sumr_149(2) or sumr_149(3) or sumr_149(4) or sumr_149(5) or sumr_149(6) or sumr_149(7) or sumr_149(8) or sumr_149(9));
E(873)<=not ( sumr_150(0) or sumr_150(1) or sumr_150(2) or sumr_150(3) or sumr_150(4) or sumr_150(5) or sumr_150(6) or sumr_150(7) or sumr_150(8) or sumr_150(9));
E(872)<=not ( sumr_151(0) or sumr_151(1) or sumr_151(2) or sumr_151(3) or sumr_151(4) or sumr_151(5) or sumr_151(6) or sumr_151(7) or sumr_151(8) or sumr_151(9));
E(871)<=not ( sumr_152(0) or sumr_152(1) or sumr_152(2) or sumr_152(3) or sumr_152(4) or sumr_152(5) or sumr_152(6) or sumr_152(7) or sumr_152(8) or sumr_152(9));
E(870)<=not ( sumr_153(0) or sumr_153(1) or sumr_153(2) or sumr_153(3) or sumr_153(4) or sumr_153(5) or sumr_153(6) or sumr_153(7) or sumr_153(8) or sumr_153(9));
E(869)<=not ( sumr_154(0) or sumr_154(1) or sumr_154(2) or sumr_154(3) or sumr_154(4) or sumr_154(5) or sumr_154(6) or sumr_154(7) or sumr_154(8) or sumr_154(9));
E(868)<=not ( sumr_155(0) or sumr_155(1) or sumr_155(2) or sumr_155(3) or sumr_155(4) or sumr_155(5) or sumr_155(6) or sumr_155(7) or sumr_155(8) or sumr_155(9));
E(867)<=not ( sumr_156(0) or sumr_156(1) or sumr_156(2) or sumr_156(3) or sumr_156(4) or sumr_156(5) or sumr_156(6) or sumr_156(7) or sumr_156(8) or sumr_156(9));
E(866)<=not ( sumr_157(0) or sumr_157(1) or sumr_157(2) or sumr_157(3) or sumr_157(4) or sumr_157(5) or sumr_157(6) or sumr_157(7) or sumr_157(8) or sumr_157(9));
E(865)<=not ( sumr_158(0) or sumr_158(1) or sumr_158(2) or sumr_158(3) or sumr_158(4) or sumr_158(5) or sumr_158(6) or sumr_158(7) or sumr_158(8) or sumr_158(9));
E(864)<=not ( sumr_159(0) or sumr_159(1) or sumr_159(2) or sumr_159(3) or sumr_159(4) or sumr_159(5) or sumr_159(6) or sumr_159(7) or sumr_159(8) or sumr_159(9));
E(863)<=not ( sumr_160(0) or sumr_160(1) or sumr_160(2) or sumr_160(3) or sumr_160(4) or sumr_160(5) or sumr_160(6) or sumr_160(7) or sumr_160(8) or sumr_160(9));
E(862)<=not ( sumr_161(0) or sumr_161(1) or sumr_161(2) or sumr_161(3) or sumr_161(4) or sumr_161(5) or sumr_161(6) or sumr_161(7) or sumr_161(8) or sumr_161(9));
E(861)<=not ( sumr_162(0) or sumr_162(1) or sumr_162(2) or sumr_162(3) or sumr_162(4) or sumr_162(5) or sumr_162(6) or sumr_162(7) or sumr_162(8) or sumr_162(9));
E(860)<=not ( sumr_163(0) or sumr_163(1) or sumr_163(2) or sumr_163(3) or sumr_163(4) or sumr_163(5) or sumr_163(6) or sumr_163(7) or sumr_163(8) or sumr_163(9));
E(859)<=not ( sumr_164(0) or sumr_164(1) or sumr_164(2) or sumr_164(3) or sumr_164(4) or sumr_164(5) or sumr_164(6) or sumr_164(7) or sumr_164(8) or sumr_164(9));
E(858)<=not ( sumr_165(0) or sumr_165(1) or sumr_165(2) or sumr_165(3) or sumr_165(4) or sumr_165(5) or sumr_165(6) or sumr_165(7) or sumr_165(8) or sumr_165(9));
E(857)<=not ( sumr_166(0) or sumr_166(1) or sumr_166(2) or sumr_166(3) or sumr_166(4) or sumr_166(5) or sumr_166(6) or sumr_166(7) or sumr_166(8) or sumr_166(9));
E(856)<=not ( sumr_167(0) or sumr_167(1) or sumr_167(2) or sumr_167(3) or sumr_167(4) or sumr_167(5) or sumr_167(6) or sumr_167(7) or sumr_167(8) or sumr_167(9));
E(855)<=not ( sumr_168(0) or sumr_168(1) or sumr_168(2) or sumr_168(3) or sumr_168(4) or sumr_168(5) or sumr_168(6) or sumr_168(7) or sumr_168(8) or sumr_168(9));
E(854)<=not ( sumr_169(0) or sumr_169(1) or sumr_169(2) or sumr_169(3) or sumr_169(4) or sumr_169(5) or sumr_169(6) or sumr_169(7) or sumr_169(8) or sumr_169(9));
E(853)<=not ( sumr_170(0) or sumr_170(1) or sumr_170(2) or sumr_170(3) or sumr_170(4) or sumr_170(5) or sumr_170(6) or sumr_170(7) or sumr_170(8) or sumr_170(9));
E(852)<=not ( sumr_171(0) or sumr_171(1) or sumr_171(2) or sumr_171(3) or sumr_171(4) or sumr_171(5) or sumr_171(6) or sumr_171(7) or sumr_171(8) or sumr_171(9));
E(851)<=not ( sumr_172(0) or sumr_172(1) or sumr_172(2) or sumr_172(3) or sumr_172(4) or sumr_172(5) or sumr_172(6) or sumr_172(7) or sumr_172(8) or sumr_172(9));
E(850)<=not ( sumr_173(0) or sumr_173(1) or sumr_173(2) or sumr_173(3) or sumr_173(4) or sumr_173(5) or sumr_173(6) or sumr_173(7) or sumr_173(8) or sumr_173(9));
E(849)<=not ( sumr_174(0) or sumr_174(1) or sumr_174(2) or sumr_174(3) or sumr_174(4) or sumr_174(5) or sumr_174(6) or sumr_174(7) or sumr_174(8) or sumr_174(9));
E(848)<=not ( sumr_175(0) or sumr_175(1) or sumr_175(2) or sumr_175(3) or sumr_175(4) or sumr_175(5) or sumr_175(6) or sumr_175(7) or sumr_175(8) or sumr_175(9));
E(847)<=not ( sumr_176(0) or sumr_176(1) or sumr_176(2) or sumr_176(3) or sumr_176(4) or sumr_176(5) or sumr_176(6) or sumr_176(7) or sumr_176(8) or sumr_176(9));
E(846)<=not ( sumr_177(0) or sumr_177(1) or sumr_177(2) or sumr_177(3) or sumr_177(4) or sumr_177(5) or sumr_177(6) or sumr_177(7) or sumr_177(8) or sumr_177(9));
E(845)<=not ( sumr_178(0) or sumr_178(1) or sumr_178(2) or sumr_178(3) or sumr_178(4) or sumr_178(5) or sumr_178(6) or sumr_178(7) or sumr_178(8) or sumr_178(9));
E(844)<=not ( sumr_179(0) or sumr_179(1) or sumr_179(2) or sumr_179(3) or sumr_179(4) or sumr_179(5) or sumr_179(6) or sumr_179(7) or sumr_179(8) or sumr_179(9));
E(843)<=not ( sumr_180(0) or sumr_180(1) or sumr_180(2) or sumr_180(3) or sumr_180(4) or sumr_180(5) or sumr_180(6) or sumr_180(7) or sumr_180(8) or sumr_180(9));
E(842)<=not ( sumr_181(0) or sumr_181(1) or sumr_181(2) or sumr_181(3) or sumr_181(4) or sumr_181(5) or sumr_181(6) or sumr_181(7) or sumr_181(8) or sumr_181(9));
E(841)<=not ( sumr_182(0) or sumr_182(1) or sumr_182(2) or sumr_182(3) or sumr_182(4) or sumr_182(5) or sumr_182(6) or sumr_182(7) or sumr_182(8) or sumr_182(9));
E(840)<=not ( sumr_183(0) or sumr_183(1) or sumr_183(2) or sumr_183(3) or sumr_183(4) or sumr_183(5) or sumr_183(6) or sumr_183(7) or sumr_183(8) or sumr_183(9));
E(839)<=not ( sumr_184(0) or sumr_184(1) or sumr_184(2) or sumr_184(3) or sumr_184(4) or sumr_184(5) or sumr_184(6) or sumr_184(7) or sumr_184(8) or sumr_184(9));
E(838)<=not ( sumr_185(0) or sumr_185(1) or sumr_185(2) or sumr_185(3) or sumr_185(4) or sumr_185(5) or sumr_185(6) or sumr_185(7) or sumr_185(8) or sumr_185(9));
E(837)<=not ( sumr_186(0) or sumr_186(1) or sumr_186(2) or sumr_186(3) or sumr_186(4) or sumr_186(5) or sumr_186(6) or sumr_186(7) or sumr_186(8) or sumr_186(9));
E(836)<=not ( sumr_187(0) or sumr_187(1) or sumr_187(2) or sumr_187(3) or sumr_187(4) or sumr_187(5) or sumr_187(6) or sumr_187(7) or sumr_187(8) or sumr_187(9));
E(835)<=not ( sumr_188(0) or sumr_188(1) or sumr_188(2) or sumr_188(3) or sumr_188(4) or sumr_188(5) or sumr_188(6) or sumr_188(7) or sumr_188(8) or sumr_188(9));
E(834)<=not ( sumr_189(0) or sumr_189(1) or sumr_189(2) or sumr_189(3) or sumr_189(4) or sumr_189(5) or sumr_189(6) or sumr_189(7) or sumr_189(8) or sumr_189(9));
E(833)<=not ( sumr_190(0) or sumr_190(1) or sumr_190(2) or sumr_190(3) or sumr_190(4) or sumr_190(5) or sumr_190(6) or sumr_190(7) or sumr_190(8) or sumr_190(9));
E(832)<=not ( sumr_191(0) or sumr_191(1) or sumr_191(2) or sumr_191(3) or sumr_191(4) or sumr_191(5) or sumr_191(6) or sumr_191(7) or sumr_191(8) or sumr_191(9));
E(831)<=not ( sumr_192(0) or sumr_192(1) or sumr_192(2) or sumr_192(3) or sumr_192(4) or sumr_192(5) or sumr_192(6) or sumr_192(7) or sumr_192(8) or sumr_192(9));
E(830)<=not ( sumr_193(0) or sumr_193(1) or sumr_193(2) or sumr_193(3) or sumr_193(4) or sumr_193(5) or sumr_193(6) or sumr_193(7) or sumr_193(8) or sumr_193(9));
E(829)<=not ( sumr_194(0) or sumr_194(1) or sumr_194(2) or sumr_194(3) or sumr_194(4) or sumr_194(5) or sumr_194(6) or sumr_194(7) or sumr_194(8) or sumr_194(9));
E(828)<=not ( sumr_195(0) or sumr_195(1) or sumr_195(2) or sumr_195(3) or sumr_195(4) or sumr_195(5) or sumr_195(6) or sumr_195(7) or sumr_195(8) or sumr_195(9));
E(827)<=not ( sumr_196(0) or sumr_196(1) or sumr_196(2) or sumr_196(3) or sumr_196(4) or sumr_196(5) or sumr_196(6) or sumr_196(7) or sumr_196(8) or sumr_196(9));
E(826)<=not ( sumr_197(0) or sumr_197(1) or sumr_197(2) or sumr_197(3) or sumr_197(4) or sumr_197(5) or sumr_197(6) or sumr_197(7) or sumr_197(8) or sumr_197(9));
E(825)<=not ( sumr_198(0) or sumr_198(1) or sumr_198(2) or sumr_198(3) or sumr_198(4) or sumr_198(5) or sumr_198(6) or sumr_198(7) or sumr_198(8) or sumr_198(9));
E(824)<=not ( sumr_199(0) or sumr_199(1) or sumr_199(2) or sumr_199(3) or sumr_199(4) or sumr_199(5) or sumr_199(6) or sumr_199(7) or sumr_199(8) or sumr_199(9));
E(823)<=not ( sumr_200(0) or sumr_200(1) or sumr_200(2) or sumr_200(3) or sumr_200(4) or sumr_200(5) or sumr_200(6) or sumr_200(7) or sumr_200(8) or sumr_200(9));
E(822)<=not ( sumr_201(0) or sumr_201(1) or sumr_201(2) or sumr_201(3) or sumr_201(4) or sumr_201(5) or sumr_201(6) or sumr_201(7) or sumr_201(8) or sumr_201(9));
E(821)<=not ( sumr_202(0) or sumr_202(1) or sumr_202(2) or sumr_202(3) or sumr_202(4) or sumr_202(5) or sumr_202(6) or sumr_202(7) or sumr_202(8) or sumr_202(9));
E(820)<=not ( sumr_203(0) or sumr_203(1) or sumr_203(2) or sumr_203(3) or sumr_203(4) or sumr_203(5) or sumr_203(6) or sumr_203(7) or sumr_203(8) or sumr_203(9));
E(819)<=not ( sumr_204(0) or sumr_204(1) or sumr_204(2) or sumr_204(3) or sumr_204(4) or sumr_204(5) or sumr_204(6) or sumr_204(7) or sumr_204(8) or sumr_204(9));
E(818)<=not ( sumr_205(0) or sumr_205(1) or sumr_205(2) or sumr_205(3) or sumr_205(4) or sumr_205(5) or sumr_205(6) or sumr_205(7) or sumr_205(8) or sumr_205(9));
E(817)<=not ( sumr_206(0) or sumr_206(1) or sumr_206(2) or sumr_206(3) or sumr_206(4) or sumr_206(5) or sumr_206(6) or sumr_206(7) or sumr_206(8) or sumr_206(9));
E(816)<=not ( sumr_207(0) or sumr_207(1) or sumr_207(2) or sumr_207(3) or sumr_207(4) or sumr_207(5) or sumr_207(6) or sumr_207(7) or sumr_207(8) or sumr_207(9));
E(815)<=not ( sumr_208(0) or sumr_208(1) or sumr_208(2) or sumr_208(3) or sumr_208(4) or sumr_208(5) or sumr_208(6) or sumr_208(7) or sumr_208(8) or sumr_208(9));
E(814)<=not ( sumr_209(0) or sumr_209(1) or sumr_209(2) or sumr_209(3) or sumr_209(4) or sumr_209(5) or sumr_209(6) or sumr_209(7) or sumr_209(8) or sumr_209(9));
E(813)<=not ( sumr_210(0) or sumr_210(1) or sumr_210(2) or sumr_210(3) or sumr_210(4) or sumr_210(5) or sumr_210(6) or sumr_210(7) or sumr_210(8) or sumr_210(9));
E(812)<=not ( sumr_211(0) or sumr_211(1) or sumr_211(2) or sumr_211(3) or sumr_211(4) or sumr_211(5) or sumr_211(6) or sumr_211(7) or sumr_211(8) or sumr_211(9));
E(811)<=not ( sumr_212(0) or sumr_212(1) or sumr_212(2) or sumr_212(3) or sumr_212(4) or sumr_212(5) or sumr_212(6) or sumr_212(7) or sumr_212(8) or sumr_212(9));
E(810)<=not ( sumr_213(0) or sumr_213(1) or sumr_213(2) or sumr_213(3) or sumr_213(4) or sumr_213(5) or sumr_213(6) or sumr_213(7) or sumr_213(8) or sumr_213(9));
E(809)<=not ( sumr_214(0) or sumr_214(1) or sumr_214(2) or sumr_214(3) or sumr_214(4) or sumr_214(5) or sumr_214(6) or sumr_214(7) or sumr_214(8) or sumr_214(9));
E(808)<=not ( sumr_215(0) or sumr_215(1) or sumr_215(2) or sumr_215(3) or sumr_215(4) or sumr_215(5) or sumr_215(6) or sumr_215(7) or sumr_215(8) or sumr_215(9));
E(807)<=not ( sumr_216(0) or sumr_216(1) or sumr_216(2) or sumr_216(3) or sumr_216(4) or sumr_216(5) or sumr_216(6) or sumr_216(7) or sumr_216(8) or sumr_216(9));
E(806)<=not ( sumr_217(0) or sumr_217(1) or sumr_217(2) or sumr_217(3) or sumr_217(4) or sumr_217(5) or sumr_217(6) or sumr_217(7) or sumr_217(8) or sumr_217(9));
E(805)<=not ( sumr_218(0) or sumr_218(1) or sumr_218(2) or sumr_218(3) or sumr_218(4) or sumr_218(5) or sumr_218(6) or sumr_218(7) or sumr_218(8) or sumr_218(9));
E(804)<=not ( sumr_219(0) or sumr_219(1) or sumr_219(2) or sumr_219(3) or sumr_219(4) or sumr_219(5) or sumr_219(6) or sumr_219(7) or sumr_219(8) or sumr_219(9));
E(803)<=not ( sumr_220(0) or sumr_220(1) or sumr_220(2) or sumr_220(3) or sumr_220(4) or sumr_220(5) or sumr_220(6) or sumr_220(7) or sumr_220(8) or sumr_220(9));
E(802)<=not ( sumr_221(0) or sumr_221(1) or sumr_221(2) or sumr_221(3) or sumr_221(4) or sumr_221(5) or sumr_221(6) or sumr_221(7) or sumr_221(8) or sumr_221(9));
E(801)<=not ( sumr_222(0) or sumr_222(1) or sumr_222(2) or sumr_222(3) or sumr_222(4) or sumr_222(5) or sumr_222(6) or sumr_222(7) or sumr_222(8) or sumr_222(9));
E(800)<=not ( sumr_223(0) or sumr_223(1) or sumr_223(2) or sumr_223(3) or sumr_223(4) or sumr_223(5) or sumr_223(6) or sumr_223(7) or sumr_223(8) or sumr_223(9));
E(799)<=not ( sumr_224(0) or sumr_224(1) or sumr_224(2) or sumr_224(3) or sumr_224(4) or sumr_224(5) or sumr_224(6) or sumr_224(7) or sumr_224(8) or sumr_224(9));
E(798)<=not ( sumr_225(0) or sumr_225(1) or sumr_225(2) or sumr_225(3) or sumr_225(4) or sumr_225(5) or sumr_225(6) or sumr_225(7) or sumr_225(8) or sumr_225(9));
E(797)<=not ( sumr_226(0) or sumr_226(1) or sumr_226(2) or sumr_226(3) or sumr_226(4) or sumr_226(5) or sumr_226(6) or sumr_226(7) or sumr_226(8) or sumr_226(9));
E(796)<=not ( sumr_227(0) or sumr_227(1) or sumr_227(2) or sumr_227(3) or sumr_227(4) or sumr_227(5) or sumr_227(6) or sumr_227(7) or sumr_227(8) or sumr_227(9));
E(795)<=not ( sumr_228(0) or sumr_228(1) or sumr_228(2) or sumr_228(3) or sumr_228(4) or sumr_228(5) or sumr_228(6) or sumr_228(7) or sumr_228(8) or sumr_228(9));
E(794)<=not ( sumr_229(0) or sumr_229(1) or sumr_229(2) or sumr_229(3) or sumr_229(4) or sumr_229(5) or sumr_229(6) or sumr_229(7) or sumr_229(8) or sumr_229(9));
E(793)<=not ( sumr_230(0) or sumr_230(1) or sumr_230(2) or sumr_230(3) or sumr_230(4) or sumr_230(5) or sumr_230(6) or sumr_230(7) or sumr_230(8) or sumr_230(9));
E(792)<=not ( sumr_231(0) or sumr_231(1) or sumr_231(2) or sumr_231(3) or sumr_231(4) or sumr_231(5) or sumr_231(6) or sumr_231(7) or sumr_231(8) or sumr_231(9));
E(791)<=not ( sumr_232(0) or sumr_232(1) or sumr_232(2) or sumr_232(3) or sumr_232(4) or sumr_232(5) or sumr_232(6) or sumr_232(7) or sumr_232(8) or sumr_232(9));
E(790)<=not ( sumr_233(0) or sumr_233(1) or sumr_233(2) or sumr_233(3) or sumr_233(4) or sumr_233(5) or sumr_233(6) or sumr_233(7) or sumr_233(8) or sumr_233(9));
E(789)<=not ( sumr_234(0) or sumr_234(1) or sumr_234(2) or sumr_234(3) or sumr_234(4) or sumr_234(5) or sumr_234(6) or sumr_234(7) or sumr_234(8) or sumr_234(9));
E(788)<=not ( sumr_235(0) or sumr_235(1) or sumr_235(2) or sumr_235(3) or sumr_235(4) or sumr_235(5) or sumr_235(6) or sumr_235(7) or sumr_235(8) or sumr_235(9));
E(787)<=not ( sumr_236(0) or sumr_236(1) or sumr_236(2) or sumr_236(3) or sumr_236(4) or sumr_236(5) or sumr_236(6) or sumr_236(7) or sumr_236(8) or sumr_236(9));
E(786)<=not ( sumr_237(0) or sumr_237(1) or sumr_237(2) or sumr_237(3) or sumr_237(4) or sumr_237(5) or sumr_237(6) or sumr_237(7) or sumr_237(8) or sumr_237(9));
E(785)<=not ( sumr_238(0) or sumr_238(1) or sumr_238(2) or sumr_238(3) or sumr_238(4) or sumr_238(5) or sumr_238(6) or sumr_238(7) or sumr_238(8) or sumr_238(9));
E(784)<=not ( sumr_239(0) or sumr_239(1) or sumr_239(2) or sumr_239(3) or sumr_239(4) or sumr_239(5) or sumr_239(6) or sumr_239(7) or sumr_239(8) or sumr_239(9));
E(783)<=not ( sumr_240(0) or sumr_240(1) or sumr_240(2) or sumr_240(3) or sumr_240(4) or sumr_240(5) or sumr_240(6) or sumr_240(7) or sumr_240(8) or sumr_240(9));
E(782)<=not ( sumr_241(0) or sumr_241(1) or sumr_241(2) or sumr_241(3) or sumr_241(4) or sumr_241(5) or sumr_241(6) or sumr_241(7) or sumr_241(8) or sumr_241(9));
E(781)<=not ( sumr_242(0) or sumr_242(1) or sumr_242(2) or sumr_242(3) or sumr_242(4) or sumr_242(5) or sumr_242(6) or sumr_242(7) or sumr_242(8) or sumr_242(9));
E(780)<=not ( sumr_243(0) or sumr_243(1) or sumr_243(2) or sumr_243(3) or sumr_243(4) or sumr_243(5) or sumr_243(6) or sumr_243(7) or sumr_243(8) or sumr_243(9));
E(779)<=not ( sumr_244(0) or sumr_244(1) or sumr_244(2) or sumr_244(3) or sumr_244(4) or sumr_244(5) or sumr_244(6) or sumr_244(7) or sumr_244(8) or sumr_244(9));
E(778)<=not ( sumr_245(0) or sumr_245(1) or sumr_245(2) or sumr_245(3) or sumr_245(4) or sumr_245(5) or sumr_245(6) or sumr_245(7) or sumr_245(8) or sumr_245(9));
E(777)<=not ( sumr_246(0) or sumr_246(1) or sumr_246(2) or sumr_246(3) or sumr_246(4) or sumr_246(5) or sumr_246(6) or sumr_246(7) or sumr_246(8) or sumr_246(9));
E(776)<=not ( sumr_247(0) or sumr_247(1) or sumr_247(2) or sumr_247(3) or sumr_247(4) or sumr_247(5) or sumr_247(6) or sumr_247(7) or sumr_247(8) or sumr_247(9));
E(775)<=not ( sumr_248(0) or sumr_248(1) or sumr_248(2) or sumr_248(3) or sumr_248(4) or sumr_248(5) or sumr_248(6) or sumr_248(7) or sumr_248(8) or sumr_248(9));
E(774)<=not ( sumr_249(0) or sumr_249(1) or sumr_249(2) or sumr_249(3) or sumr_249(4) or sumr_249(5) or sumr_249(6) or sumr_249(7) or sumr_249(8) or sumr_249(9));
E(773)<=not ( sumr_250(0) or sumr_250(1) or sumr_250(2) or sumr_250(3) or sumr_250(4) or sumr_250(5) or sumr_250(6) or sumr_250(7) or sumr_250(8) or sumr_250(9));
E(772)<=not ( sumr_251(0) or sumr_251(1) or sumr_251(2) or sumr_251(3) or sumr_251(4) or sumr_251(5) or sumr_251(6) or sumr_251(7) or sumr_251(8) or sumr_251(9));
E(771)<=not ( sumr_252(0) or sumr_252(1) or sumr_252(2) or sumr_252(3) or sumr_252(4) or sumr_252(5) or sumr_252(6) or sumr_252(7) or sumr_252(8) or sumr_252(9));
E(770)<=not ( sumr_253(0) or sumr_253(1) or sumr_253(2) or sumr_253(3) or sumr_253(4) or sumr_253(5) or sumr_253(6) or sumr_253(7) or sumr_253(8) or sumr_253(9));
E(769)<=not ( sumr_254(0) or sumr_254(1) or sumr_254(2) or sumr_254(3) or sumr_254(4) or sumr_254(5) or sumr_254(6) or sumr_254(7) or sumr_254(8) or sumr_254(9));
E(768)<=not ( sumr_255(0) or sumr_255(1) or sumr_255(2) or sumr_255(3) or sumr_255(4) or sumr_255(5) or sumr_255(6) or sumr_255(7) or sumr_255(8) or sumr_255(9));
E(767)<=not ( sumr_256(0) or sumr_256(1) or sumr_256(2) or sumr_256(3) or sumr_256(4) or sumr_256(5) or sumr_256(6) or sumr_256(7) or sumr_256(8) or sumr_256(9));
E(766)<=not ( sumr_257(0) or sumr_257(1) or sumr_257(2) or sumr_257(3) or sumr_257(4) or sumr_257(5) or sumr_257(6) or sumr_257(7) or sumr_257(8) or sumr_257(9));
E(765)<=not ( sumr_258(0) or sumr_258(1) or sumr_258(2) or sumr_258(3) or sumr_258(4) or sumr_258(5) or sumr_258(6) or sumr_258(7) or sumr_258(8) or sumr_258(9));
E(764)<=not ( sumr_259(0) or sumr_259(1) or sumr_259(2) or sumr_259(3) or sumr_259(4) or sumr_259(5) or sumr_259(6) or sumr_259(7) or sumr_259(8) or sumr_259(9));
E(763)<=not ( sumr_260(0) or sumr_260(1) or sumr_260(2) or sumr_260(3) or sumr_260(4) or sumr_260(5) or sumr_260(6) or sumr_260(7) or sumr_260(8) or sumr_260(9));
E(762)<=not ( sumr_261(0) or sumr_261(1) or sumr_261(2) or sumr_261(3) or sumr_261(4) or sumr_261(5) or sumr_261(6) or sumr_261(7) or sumr_261(8) or sumr_261(9));
E(761)<=not ( sumr_262(0) or sumr_262(1) or sumr_262(2) or sumr_262(3) or sumr_262(4) or sumr_262(5) or sumr_262(6) or sumr_262(7) or sumr_262(8) or sumr_262(9));
E(760)<=not ( sumr_263(0) or sumr_263(1) or sumr_263(2) or sumr_263(3) or sumr_263(4) or sumr_263(5) or sumr_263(6) or sumr_263(7) or sumr_263(8) or sumr_263(9));
E(759)<=not ( sumr_264(0) or sumr_264(1) or sumr_264(2) or sumr_264(3) or sumr_264(4) or sumr_264(5) or sumr_264(6) or sumr_264(7) or sumr_264(8) or sumr_264(9));
E(758)<=not ( sumr_265(0) or sumr_265(1) or sumr_265(2) or sumr_265(3) or sumr_265(4) or sumr_265(5) or sumr_265(6) or sumr_265(7) or sumr_265(8) or sumr_265(9));
E(757)<=not ( sumr_266(0) or sumr_266(1) or sumr_266(2) or sumr_266(3) or sumr_266(4) or sumr_266(5) or sumr_266(6) or sumr_266(7) or sumr_266(8) or sumr_266(9));
E(756)<=not ( sumr_267(0) or sumr_267(1) or sumr_267(2) or sumr_267(3) or sumr_267(4) or sumr_267(5) or sumr_267(6) or sumr_267(7) or sumr_267(8) or sumr_267(9));
E(755)<=not ( sumr_268(0) or sumr_268(1) or sumr_268(2) or sumr_268(3) or sumr_268(4) or sumr_268(5) or sumr_268(6) or sumr_268(7) or sumr_268(8) or sumr_268(9));
E(754)<=not ( sumr_269(0) or sumr_269(1) or sumr_269(2) or sumr_269(3) or sumr_269(4) or sumr_269(5) or sumr_269(6) or sumr_269(7) or sumr_269(8) or sumr_269(9));
E(753)<=not ( sumr_270(0) or sumr_270(1) or sumr_270(2) or sumr_270(3) or sumr_270(4) or sumr_270(5) or sumr_270(6) or sumr_270(7) or sumr_270(8) or sumr_270(9));
E(752)<=not ( sumr_271(0) or sumr_271(1) or sumr_271(2) or sumr_271(3) or sumr_271(4) or sumr_271(5) or sumr_271(6) or sumr_271(7) or sumr_271(8) or sumr_271(9));
E(751)<=not ( sumr_272(0) or sumr_272(1) or sumr_272(2) or sumr_272(3) or sumr_272(4) or sumr_272(5) or sumr_272(6) or sumr_272(7) or sumr_272(8) or sumr_272(9));
E(750)<=not ( sumr_273(0) or sumr_273(1) or sumr_273(2) or sumr_273(3) or sumr_273(4) or sumr_273(5) or sumr_273(6) or sumr_273(7) or sumr_273(8) or sumr_273(9));
E(749)<=not ( sumr_274(0) or sumr_274(1) or sumr_274(2) or sumr_274(3) or sumr_274(4) or sumr_274(5) or sumr_274(6) or sumr_274(7) or sumr_274(8) or sumr_274(9));
E(748)<=not ( sumr_275(0) or sumr_275(1) or sumr_275(2) or sumr_275(3) or sumr_275(4) or sumr_275(5) or sumr_275(6) or sumr_275(7) or sumr_275(8) or sumr_275(9));
E(747)<=not ( sumr_276(0) or sumr_276(1) or sumr_276(2) or sumr_276(3) or sumr_276(4) or sumr_276(5) or sumr_276(6) or sumr_276(7) or sumr_276(8) or sumr_276(9));
E(746)<=not ( sumr_277(0) or sumr_277(1) or sumr_277(2) or sumr_277(3) or sumr_277(4) or sumr_277(5) or sumr_277(6) or sumr_277(7) or sumr_277(8) or sumr_277(9));
E(745)<=not ( sumr_278(0) or sumr_278(1) or sumr_278(2) or sumr_278(3) or sumr_278(4) or sumr_278(5) or sumr_278(6) or sumr_278(7) or sumr_278(8) or sumr_278(9));
E(744)<=not ( sumr_279(0) or sumr_279(1) or sumr_279(2) or sumr_279(3) or sumr_279(4) or sumr_279(5) or sumr_279(6) or sumr_279(7) or sumr_279(8) or sumr_279(9));
E(743)<=not ( sumr_280(0) or sumr_280(1) or sumr_280(2) or sumr_280(3) or sumr_280(4) or sumr_280(5) or sumr_280(6) or sumr_280(7) or sumr_280(8) or sumr_280(9));
E(742)<=not ( sumr_281(0) or sumr_281(1) or sumr_281(2) or sumr_281(3) or sumr_281(4) or sumr_281(5) or sumr_281(6) or sumr_281(7) or sumr_281(8) or sumr_281(9));
E(741)<=not ( sumr_282(0) or sumr_282(1) or sumr_282(2) or sumr_282(3) or sumr_282(4) or sumr_282(5) or sumr_282(6) or sumr_282(7) or sumr_282(8) or sumr_282(9));
E(740)<=not ( sumr_283(0) or sumr_283(1) or sumr_283(2) or sumr_283(3) or sumr_283(4) or sumr_283(5) or sumr_283(6) or sumr_283(7) or sumr_283(8) or sumr_283(9));
E(739)<=not ( sumr_284(0) or sumr_284(1) or sumr_284(2) or sumr_284(3) or sumr_284(4) or sumr_284(5) or sumr_284(6) or sumr_284(7) or sumr_284(8) or sumr_284(9));
E(738)<=not ( sumr_285(0) or sumr_285(1) or sumr_285(2) or sumr_285(3) or sumr_285(4) or sumr_285(5) or sumr_285(6) or sumr_285(7) or sumr_285(8) or sumr_285(9));
E(737)<=not ( sumr_286(0) or sumr_286(1) or sumr_286(2) or sumr_286(3) or sumr_286(4) or sumr_286(5) or sumr_286(6) or sumr_286(7) or sumr_286(8) or sumr_286(9));
E(736)<=not ( sumr_287(0) or sumr_287(1) or sumr_287(2) or sumr_287(3) or sumr_287(4) or sumr_287(5) or sumr_287(6) or sumr_287(7) or sumr_287(8) or sumr_287(9));
E(735)<=not ( sumr_288(0) or sumr_288(1) or sumr_288(2) or sumr_288(3) or sumr_288(4) or sumr_288(5) or sumr_288(6) or sumr_288(7) or sumr_288(8) or sumr_288(9));
E(734)<=not ( sumr_289(0) or sumr_289(1) or sumr_289(2) or sumr_289(3) or sumr_289(4) or sumr_289(5) or sumr_289(6) or sumr_289(7) or sumr_289(8) or sumr_289(9));
E(733)<=not ( sumr_290(0) or sumr_290(1) or sumr_290(2) or sumr_290(3) or sumr_290(4) or sumr_290(5) or sumr_290(6) or sumr_290(7) or sumr_290(8) or sumr_290(9));
E(732)<=not ( sumr_291(0) or sumr_291(1) or sumr_291(2) or sumr_291(3) or sumr_291(4) or sumr_291(5) or sumr_291(6) or sumr_291(7) or sumr_291(8) or sumr_291(9));
E(731)<=not ( sumr_292(0) or sumr_292(1) or sumr_292(2) or sumr_292(3) or sumr_292(4) or sumr_292(5) or sumr_292(6) or sumr_292(7) or sumr_292(8) or sumr_292(9));
E(730)<=not ( sumr_293(0) or sumr_293(1) or sumr_293(2) or sumr_293(3) or sumr_293(4) or sumr_293(5) or sumr_293(6) or sumr_293(7) or sumr_293(8) or sumr_293(9));
E(729)<=not ( sumr_294(0) or sumr_294(1) or sumr_294(2) or sumr_294(3) or sumr_294(4) or sumr_294(5) or sumr_294(6) or sumr_294(7) or sumr_294(8) or sumr_294(9));
E(728)<=not ( sumr_295(0) or sumr_295(1) or sumr_295(2) or sumr_295(3) or sumr_295(4) or sumr_295(5) or sumr_295(6) or sumr_295(7) or sumr_295(8) or sumr_295(9));
E(727)<=not ( sumr_296(0) or sumr_296(1) or sumr_296(2) or sumr_296(3) or sumr_296(4) or sumr_296(5) or sumr_296(6) or sumr_296(7) or sumr_296(8) or sumr_296(9));
E(726)<=not ( sumr_297(0) or sumr_297(1) or sumr_297(2) or sumr_297(3) or sumr_297(4) or sumr_297(5) or sumr_297(6) or sumr_297(7) or sumr_297(8) or sumr_297(9));
E(725)<=not ( sumr_298(0) or sumr_298(1) or sumr_298(2) or sumr_298(3) or sumr_298(4) or sumr_298(5) or sumr_298(6) or sumr_298(7) or sumr_298(8) or sumr_298(9));
E(724)<=not ( sumr_299(0) or sumr_299(1) or sumr_299(2) or sumr_299(3) or sumr_299(4) or sumr_299(5) or sumr_299(6) or sumr_299(7) or sumr_299(8) or sumr_299(9));
E(723)<=not ( sumr_300(0) or sumr_300(1) or sumr_300(2) or sumr_300(3) or sumr_300(4) or sumr_300(5) or sumr_300(6) or sumr_300(7) or sumr_300(8) or sumr_300(9));
E(722)<=not ( sumr_301(0) or sumr_301(1) or sumr_301(2) or sumr_301(3) or sumr_301(4) or sumr_301(5) or sumr_301(6) or sumr_301(7) or sumr_301(8) or sumr_301(9));
E(721)<=not ( sumr_302(0) or sumr_302(1) or sumr_302(2) or sumr_302(3) or sumr_302(4) or sumr_302(5) or sumr_302(6) or sumr_302(7) or sumr_302(8) or sumr_302(9));
E(720)<=not ( sumr_303(0) or sumr_303(1) or sumr_303(2) or sumr_303(3) or sumr_303(4) or sumr_303(5) or sumr_303(6) or sumr_303(7) or sumr_303(8) or sumr_303(9));
E(719)<=not ( sumr_304(0) or sumr_304(1) or sumr_304(2) or sumr_304(3) or sumr_304(4) or sumr_304(5) or sumr_304(6) or sumr_304(7) or sumr_304(8) or sumr_304(9));
E(718)<=not ( sumr_305(0) or sumr_305(1) or sumr_305(2) or sumr_305(3) or sumr_305(4) or sumr_305(5) or sumr_305(6) or sumr_305(7) or sumr_305(8) or sumr_305(9));
E(717)<=not ( sumr_306(0) or sumr_306(1) or sumr_306(2) or sumr_306(3) or sumr_306(4) or sumr_306(5) or sumr_306(6) or sumr_306(7) or sumr_306(8) or sumr_306(9));
E(716)<=not ( sumr_307(0) or sumr_307(1) or sumr_307(2) or sumr_307(3) or sumr_307(4) or sumr_307(5) or sumr_307(6) or sumr_307(7) or sumr_307(8) or sumr_307(9));
E(715)<=not ( sumr_308(0) or sumr_308(1) or sumr_308(2) or sumr_308(3) or sumr_308(4) or sumr_308(5) or sumr_308(6) or sumr_308(7) or sumr_308(8) or sumr_308(9));
E(714)<=not ( sumr_309(0) or sumr_309(1) or sumr_309(2) or sumr_309(3) or sumr_309(4) or sumr_309(5) or sumr_309(6) or sumr_309(7) or sumr_309(8) or sumr_309(9));
E(713)<=not ( sumr_310(0) or sumr_310(1) or sumr_310(2) or sumr_310(3) or sumr_310(4) or sumr_310(5) or sumr_310(6) or sumr_310(7) or sumr_310(8) or sumr_310(9));
E(712)<=not ( sumr_311(0) or sumr_311(1) or sumr_311(2) or sumr_311(3) or sumr_311(4) or sumr_311(5) or sumr_311(6) or sumr_311(7) or sumr_311(8) or sumr_311(9));
E(711)<=not ( sumr_312(0) or sumr_312(1) or sumr_312(2) or sumr_312(3) or sumr_312(4) or sumr_312(5) or sumr_312(6) or sumr_312(7) or sumr_312(8) or sumr_312(9));
E(710)<=not ( sumr_313(0) or sumr_313(1) or sumr_313(2) or sumr_313(3) or sumr_313(4) or sumr_313(5) or sumr_313(6) or sumr_313(7) or sumr_313(8) or sumr_313(9));
E(709)<=not ( sumr_314(0) or sumr_314(1) or sumr_314(2) or sumr_314(3) or sumr_314(4) or sumr_314(5) or sumr_314(6) or sumr_314(7) or sumr_314(8) or sumr_314(9));
E(708)<=not ( sumr_315(0) or sumr_315(1) or sumr_315(2) or sumr_315(3) or sumr_315(4) or sumr_315(5) or sumr_315(6) or sumr_315(7) or sumr_315(8) or sumr_315(9));
E(707)<=not ( sumr_316(0) or sumr_316(1) or sumr_316(2) or sumr_316(3) or sumr_316(4) or sumr_316(5) or sumr_316(6) or sumr_316(7) or sumr_316(8) or sumr_316(9));
E(706)<=not ( sumr_317(0) or sumr_317(1) or sumr_317(2) or sumr_317(3) or sumr_317(4) or sumr_317(5) or sumr_317(6) or sumr_317(7) or sumr_317(8) or sumr_317(9));
E(705)<=not ( sumr_318(0) or sumr_318(1) or sumr_318(2) or sumr_318(3) or sumr_318(4) or sumr_318(5) or sumr_318(6) or sumr_318(7) or sumr_318(8) or sumr_318(9));
E(704)<=not ( sumr_319(0) or sumr_319(1) or sumr_319(2) or sumr_319(3) or sumr_319(4) or sumr_319(5) or sumr_319(6) or sumr_319(7) or sumr_319(8) or sumr_319(9));
E(703)<=not ( sumr_320(0) or sumr_320(1) or sumr_320(2) or sumr_320(3) or sumr_320(4) or sumr_320(5) or sumr_320(6) or sumr_320(7) or sumr_320(8) or sumr_320(9));
E(702)<=not ( sumr_321(0) or sumr_321(1) or sumr_321(2) or sumr_321(3) or sumr_321(4) or sumr_321(5) or sumr_321(6) or sumr_321(7) or sumr_321(8) or sumr_321(9));
E(701)<=not ( sumr_322(0) or sumr_322(1) or sumr_322(2) or sumr_322(3) or sumr_322(4) or sumr_322(5) or sumr_322(6) or sumr_322(7) or sumr_322(8) or sumr_322(9));
E(700)<=not ( sumr_323(0) or sumr_323(1) or sumr_323(2) or sumr_323(3) or sumr_323(4) or sumr_323(5) or sumr_323(6) or sumr_323(7) or sumr_323(8) or sumr_323(9));
E(699)<=not ( sumr_324(0) or sumr_324(1) or sumr_324(2) or sumr_324(3) or sumr_324(4) or sumr_324(5) or sumr_324(6) or sumr_324(7) or sumr_324(8) or sumr_324(9));
E(698)<=not ( sumr_325(0) or sumr_325(1) or sumr_325(2) or sumr_325(3) or sumr_325(4) or sumr_325(5) or sumr_325(6) or sumr_325(7) or sumr_325(8) or sumr_325(9));
E(697)<=not ( sumr_326(0) or sumr_326(1) or sumr_326(2) or sumr_326(3) or sumr_326(4) or sumr_326(5) or sumr_326(6) or sumr_326(7) or sumr_326(8) or sumr_326(9));
E(696)<=not ( sumr_327(0) or sumr_327(1) or sumr_327(2) or sumr_327(3) or sumr_327(4) or sumr_327(5) or sumr_327(6) or sumr_327(7) or sumr_327(8) or sumr_327(9));
E(695)<=not ( sumr_328(0) or sumr_328(1) or sumr_328(2) or sumr_328(3) or sumr_328(4) or sumr_328(5) or sumr_328(6) or sumr_328(7) or sumr_328(8) or sumr_328(9));
E(694)<=not ( sumr_329(0) or sumr_329(1) or sumr_329(2) or sumr_329(3) or sumr_329(4) or sumr_329(5) or sumr_329(6) or sumr_329(7) or sumr_329(8) or sumr_329(9));
E(693)<=not ( sumr_330(0) or sumr_330(1) or sumr_330(2) or sumr_330(3) or sumr_330(4) or sumr_330(5) or sumr_330(6) or sumr_330(7) or sumr_330(8) or sumr_330(9));
E(692)<=not ( sumr_331(0) or sumr_331(1) or sumr_331(2) or sumr_331(3) or sumr_331(4) or sumr_331(5) or sumr_331(6) or sumr_331(7) or sumr_331(8) or sumr_331(9));
E(691)<=not ( sumr_332(0) or sumr_332(1) or sumr_332(2) or sumr_332(3) or sumr_332(4) or sumr_332(5) or sumr_332(6) or sumr_332(7) or sumr_332(8) or sumr_332(9));
E(690)<=not ( sumr_333(0) or sumr_333(1) or sumr_333(2) or sumr_333(3) or sumr_333(4) or sumr_333(5) or sumr_333(6) or sumr_333(7) or sumr_333(8) or sumr_333(9));
E(689)<=not ( sumr_334(0) or sumr_334(1) or sumr_334(2) or sumr_334(3) or sumr_334(4) or sumr_334(5) or sumr_334(6) or sumr_334(7) or sumr_334(8) or sumr_334(9));
E(688)<=not ( sumr_335(0) or sumr_335(1) or sumr_335(2) or sumr_335(3) or sumr_335(4) or sumr_335(5) or sumr_335(6) or sumr_335(7) or sumr_335(8) or sumr_335(9));
E(687)<=not ( sumr_336(0) or sumr_336(1) or sumr_336(2) or sumr_336(3) or sumr_336(4) or sumr_336(5) or sumr_336(6) or sumr_336(7) or sumr_336(8) or sumr_336(9));
E(686)<=not ( sumr_337(0) or sumr_337(1) or sumr_337(2) or sumr_337(3) or sumr_337(4) or sumr_337(5) or sumr_337(6) or sumr_337(7) or sumr_337(8) or sumr_337(9));
E(685)<=not ( sumr_338(0) or sumr_338(1) or sumr_338(2) or sumr_338(3) or sumr_338(4) or sumr_338(5) or sumr_338(6) or sumr_338(7) or sumr_338(8) or sumr_338(9));
E(684)<=not ( sumr_339(0) or sumr_339(1) or sumr_339(2) or sumr_339(3) or sumr_339(4) or sumr_339(5) or sumr_339(6) or sumr_339(7) or sumr_339(8) or sumr_339(9));
E(683)<=not ( sumr_340(0) or sumr_340(1) or sumr_340(2) or sumr_340(3) or sumr_340(4) or sumr_340(5) or sumr_340(6) or sumr_340(7) or sumr_340(8) or sumr_340(9));
E(682)<=not ( sumr_341(0) or sumr_341(1) or sumr_341(2) or sumr_341(3) or sumr_341(4) or sumr_341(5) or sumr_341(6) or sumr_341(7) or sumr_341(8) or sumr_341(9));
E(681)<=not ( sumr_342(0) or sumr_342(1) or sumr_342(2) or sumr_342(3) or sumr_342(4) or sumr_342(5) or sumr_342(6) or sumr_342(7) or sumr_342(8) or sumr_342(9));
E(680)<=not ( sumr_343(0) or sumr_343(1) or sumr_343(2) or sumr_343(3) or sumr_343(4) or sumr_343(5) or sumr_343(6) or sumr_343(7) or sumr_343(8) or sumr_343(9));
E(679)<=not ( sumr_344(0) or sumr_344(1) or sumr_344(2) or sumr_344(3) or sumr_344(4) or sumr_344(5) or sumr_344(6) or sumr_344(7) or sumr_344(8) or sumr_344(9));
E(678)<=not ( sumr_345(0) or sumr_345(1) or sumr_345(2) or sumr_345(3) or sumr_345(4) or sumr_345(5) or sumr_345(6) or sumr_345(7) or sumr_345(8) or sumr_345(9));
E(677)<=not ( sumr_346(0) or sumr_346(1) or sumr_346(2) or sumr_346(3) or sumr_346(4) or sumr_346(5) or sumr_346(6) or sumr_346(7) or sumr_346(8) or sumr_346(9));
E(676)<=not ( sumr_347(0) or sumr_347(1) or sumr_347(2) or sumr_347(3) or sumr_347(4) or sumr_347(5) or sumr_347(6) or sumr_347(7) or sumr_347(8) or sumr_347(9));
E(675)<=not ( sumr_348(0) or sumr_348(1) or sumr_348(2) or sumr_348(3) or sumr_348(4) or sumr_348(5) or sumr_348(6) or sumr_348(7) or sumr_348(8) or sumr_348(9));
E(674)<=not ( sumr_349(0) or sumr_349(1) or sumr_349(2) or sumr_349(3) or sumr_349(4) or sumr_349(5) or sumr_349(6) or sumr_349(7) or sumr_349(8) or sumr_349(9));
E(673)<=not ( sumr_350(0) or sumr_350(1) or sumr_350(2) or sumr_350(3) or sumr_350(4) or sumr_350(5) or sumr_350(6) or sumr_350(7) or sumr_350(8) or sumr_350(9));
E(672)<=not ( sumr_351(0) or sumr_351(1) or sumr_351(2) or sumr_351(3) or sumr_351(4) or sumr_351(5) or sumr_351(6) or sumr_351(7) or sumr_351(8) or sumr_351(9));
E(671)<=not ( sumr_352(0) or sumr_352(1) or sumr_352(2) or sumr_352(3) or sumr_352(4) or sumr_352(5) or sumr_352(6) or sumr_352(7) or sumr_352(8) or sumr_352(9));
E(670)<=not ( sumr_353(0) or sumr_353(1) or sumr_353(2) or sumr_353(3) or sumr_353(4) or sumr_353(5) or sumr_353(6) or sumr_353(7) or sumr_353(8) or sumr_353(9));
E(669)<=not ( sumr_354(0) or sumr_354(1) or sumr_354(2) or sumr_354(3) or sumr_354(4) or sumr_354(5) or sumr_354(6) or sumr_354(7) or sumr_354(8) or sumr_354(9));
E(668)<=not ( sumr_355(0) or sumr_355(1) or sumr_355(2) or sumr_355(3) or sumr_355(4) or sumr_355(5) or sumr_355(6) or sumr_355(7) or sumr_355(8) or sumr_355(9));
E(667)<=not ( sumr_356(0) or sumr_356(1) or sumr_356(2) or sumr_356(3) or sumr_356(4) or sumr_356(5) or sumr_356(6) or sumr_356(7) or sumr_356(8) or sumr_356(9));
E(666)<=not ( sumr_357(0) or sumr_357(1) or sumr_357(2) or sumr_357(3) or sumr_357(4) or sumr_357(5) or sumr_357(6) or sumr_357(7) or sumr_357(8) or sumr_357(9));
E(665)<=not ( sumr_358(0) or sumr_358(1) or sumr_358(2) or sumr_358(3) or sumr_358(4) or sumr_358(5) or sumr_358(6) or sumr_358(7) or sumr_358(8) or sumr_358(9));
E(664)<=not ( sumr_359(0) or sumr_359(1) or sumr_359(2) or sumr_359(3) or sumr_359(4) or sumr_359(5) or sumr_359(6) or sumr_359(7) or sumr_359(8) or sumr_359(9));
E(663)<=not ( sumr_360(0) or sumr_360(1) or sumr_360(2) or sumr_360(3) or sumr_360(4) or sumr_360(5) or sumr_360(6) or sumr_360(7) or sumr_360(8) or sumr_360(9));
E(662)<=not ( sumr_361(0) or sumr_361(1) or sumr_361(2) or sumr_361(3) or sumr_361(4) or sumr_361(5) or sumr_361(6) or sumr_361(7) or sumr_361(8) or sumr_361(9));
E(661)<=not ( sumr_362(0) or sumr_362(1) or sumr_362(2) or sumr_362(3) or sumr_362(4) or sumr_362(5) or sumr_362(6) or sumr_362(7) or sumr_362(8) or sumr_362(9));
E(660)<=not ( sumr_363(0) or sumr_363(1) or sumr_363(2) or sumr_363(3) or sumr_363(4) or sumr_363(5) or sumr_363(6) or sumr_363(7) or sumr_363(8) or sumr_363(9));
E(659)<=not ( sumr_364(0) or sumr_364(1) or sumr_364(2) or sumr_364(3) or sumr_364(4) or sumr_364(5) or sumr_364(6) or sumr_364(7) or sumr_364(8) or sumr_364(9));
E(658)<=not ( sumr_365(0) or sumr_365(1) or sumr_365(2) or sumr_365(3) or sumr_365(4) or sumr_365(5) or sumr_365(6) or sumr_365(7) or sumr_365(8) or sumr_365(9));
E(657)<=not ( sumr_366(0) or sumr_366(1) or sumr_366(2) or sumr_366(3) or sumr_366(4) or sumr_366(5) or sumr_366(6) or sumr_366(7) or sumr_366(8) or sumr_366(9));
E(656)<=not ( sumr_367(0) or sumr_367(1) or sumr_367(2) or sumr_367(3) or sumr_367(4) or sumr_367(5) or sumr_367(6) or sumr_367(7) or sumr_367(8) or sumr_367(9));
E(655)<=not ( sumr_368(0) or sumr_368(1) or sumr_368(2) or sumr_368(3) or sumr_368(4) or sumr_368(5) or sumr_368(6) or sumr_368(7) or sumr_368(8) or sumr_368(9));
E(654)<=not ( sumr_369(0) or sumr_369(1) or sumr_369(2) or sumr_369(3) or sumr_369(4) or sumr_369(5) or sumr_369(6) or sumr_369(7) or sumr_369(8) or sumr_369(9));
E(653)<=not ( sumr_370(0) or sumr_370(1) or sumr_370(2) or sumr_370(3) or sumr_370(4) or sumr_370(5) or sumr_370(6) or sumr_370(7) or sumr_370(8) or sumr_370(9));
E(652)<=not ( sumr_371(0) or sumr_371(1) or sumr_371(2) or sumr_371(3) or sumr_371(4) or sumr_371(5) or sumr_371(6) or sumr_371(7) or sumr_371(8) or sumr_371(9));
E(651)<=not ( sumr_372(0) or sumr_372(1) or sumr_372(2) or sumr_372(3) or sumr_372(4) or sumr_372(5) or sumr_372(6) or sumr_372(7) or sumr_372(8) or sumr_372(9));
E(650)<=not ( sumr_373(0) or sumr_373(1) or sumr_373(2) or sumr_373(3) or sumr_373(4) or sumr_373(5) or sumr_373(6) or sumr_373(7) or sumr_373(8) or sumr_373(9));
E(649)<=not ( sumr_374(0) or sumr_374(1) or sumr_374(2) or sumr_374(3) or sumr_374(4) or sumr_374(5) or sumr_374(6) or sumr_374(7) or sumr_374(8) or sumr_374(9));
E(648)<=not ( sumr_375(0) or sumr_375(1) or sumr_375(2) or sumr_375(3) or sumr_375(4) or sumr_375(5) or sumr_375(6) or sumr_375(7) or sumr_375(8) or sumr_375(9));
E(647)<=not ( sumr_376(0) or sumr_376(1) or sumr_376(2) or sumr_376(3) or sumr_376(4) or sumr_376(5) or sumr_376(6) or sumr_376(7) or sumr_376(8) or sumr_376(9));
E(646)<=not ( sumr_377(0) or sumr_377(1) or sumr_377(2) or sumr_377(3) or sumr_377(4) or sumr_377(5) or sumr_377(6) or sumr_377(7) or sumr_377(8) or sumr_377(9));
E(645)<=not ( sumr_378(0) or sumr_378(1) or sumr_378(2) or sumr_378(3) or sumr_378(4) or sumr_378(5) or sumr_378(6) or sumr_378(7) or sumr_378(8) or sumr_378(9));
E(644)<=not ( sumr_379(0) or sumr_379(1) or sumr_379(2) or sumr_379(3) or sumr_379(4) or sumr_379(5) or sumr_379(6) or sumr_379(7) or sumr_379(8) or sumr_379(9));
E(643)<=not ( sumr_380(0) or sumr_380(1) or sumr_380(2) or sumr_380(3) or sumr_380(4) or sumr_380(5) or sumr_380(6) or sumr_380(7) or sumr_380(8) or sumr_380(9));
E(642)<=not ( sumr_381(0) or sumr_381(1) or sumr_381(2) or sumr_381(3) or sumr_381(4) or sumr_381(5) or sumr_381(6) or sumr_381(7) or sumr_381(8) or sumr_381(9));
E(641)<=not ( sumr_382(0) or sumr_382(1) or sumr_382(2) or sumr_382(3) or sumr_382(4) or sumr_382(5) or sumr_382(6) or sumr_382(7) or sumr_382(8) or sumr_382(9));
E(640)<=not ( sumr_383(0) or sumr_383(1) or sumr_383(2) or sumr_383(3) or sumr_383(4) or sumr_383(5) or sumr_383(6) or sumr_383(7) or sumr_383(8) or sumr_383(9));
E(639)<=not ( sumr_384(0) or sumr_384(1) or sumr_384(2) or sumr_384(3) or sumr_384(4) or sumr_384(5) or sumr_384(6) or sumr_384(7) or sumr_384(8) or sumr_384(9));
E(638)<=not ( sumr_385(0) or sumr_385(1) or sumr_385(2) or sumr_385(3) or sumr_385(4) or sumr_385(5) or sumr_385(6) or sumr_385(7) or sumr_385(8) or sumr_385(9));
E(637)<=not ( sumr_386(0) or sumr_386(1) or sumr_386(2) or sumr_386(3) or sumr_386(4) or sumr_386(5) or sumr_386(6) or sumr_386(7) or sumr_386(8) or sumr_386(9));
E(636)<=not ( sumr_387(0) or sumr_387(1) or sumr_387(2) or sumr_387(3) or sumr_387(4) or sumr_387(5) or sumr_387(6) or sumr_387(7) or sumr_387(8) or sumr_387(9));
E(635)<=not ( sumr_388(0) or sumr_388(1) or sumr_388(2) or sumr_388(3) or sumr_388(4) or sumr_388(5) or sumr_388(6) or sumr_388(7) or sumr_388(8) or sumr_388(9));
E(634)<=not ( sumr_389(0) or sumr_389(1) or sumr_389(2) or sumr_389(3) or sumr_389(4) or sumr_389(5) or sumr_389(6) or sumr_389(7) or sumr_389(8) or sumr_389(9));
E(633)<=not ( sumr_390(0) or sumr_390(1) or sumr_390(2) or sumr_390(3) or sumr_390(4) or sumr_390(5) or sumr_390(6) or sumr_390(7) or sumr_390(8) or sumr_390(9));
E(632)<=not ( sumr_391(0) or sumr_391(1) or sumr_391(2) or sumr_391(3) or sumr_391(4) or sumr_391(5) or sumr_391(6) or sumr_391(7) or sumr_391(8) or sumr_391(9));
E(631)<=not ( sumr_392(0) or sumr_392(1) or sumr_392(2) or sumr_392(3) or sumr_392(4) or sumr_392(5) or sumr_392(6) or sumr_392(7) or sumr_392(8) or sumr_392(9));
E(630)<=not ( sumr_393(0) or sumr_393(1) or sumr_393(2) or sumr_393(3) or sumr_393(4) or sumr_393(5) or sumr_393(6) or sumr_393(7) or sumr_393(8) or sumr_393(9));
E(629)<=not ( sumr_394(0) or sumr_394(1) or sumr_394(2) or sumr_394(3) or sumr_394(4) or sumr_394(5) or sumr_394(6) or sumr_394(7) or sumr_394(8) or sumr_394(9));
E(628)<=not ( sumr_395(0) or sumr_395(1) or sumr_395(2) or sumr_395(3) or sumr_395(4) or sumr_395(5) or sumr_395(6) or sumr_395(7) or sumr_395(8) or sumr_395(9));
E(627)<=not ( sumr_396(0) or sumr_396(1) or sumr_396(2) or sumr_396(3) or sumr_396(4) or sumr_396(5) or sumr_396(6) or sumr_396(7) or sumr_396(8) or sumr_396(9));
E(626)<=not ( sumr_397(0) or sumr_397(1) or sumr_397(2) or sumr_397(3) or sumr_397(4) or sumr_397(5) or sumr_397(6) or sumr_397(7) or sumr_397(8) or sumr_397(9));
E(625)<=not ( sumr_398(0) or sumr_398(1) or sumr_398(2) or sumr_398(3) or sumr_398(4) or sumr_398(5) or sumr_398(6) or sumr_398(7) or sumr_398(8) or sumr_398(9));
E(624)<=not ( sumr_399(0) or sumr_399(1) or sumr_399(2) or sumr_399(3) or sumr_399(4) or sumr_399(5) or sumr_399(6) or sumr_399(7) or sumr_399(8) or sumr_399(9));
E(623)<=not ( sumr_400(0) or sumr_400(1) or sumr_400(2) or sumr_400(3) or sumr_400(4) or sumr_400(5) or sumr_400(6) or sumr_400(7) or sumr_400(8) or sumr_400(9));
E(622)<=not ( sumr_401(0) or sumr_401(1) or sumr_401(2) or sumr_401(3) or sumr_401(4) or sumr_401(5) or sumr_401(6) or sumr_401(7) or sumr_401(8) or sumr_401(9));
E(621)<=not ( sumr_402(0) or sumr_402(1) or sumr_402(2) or sumr_402(3) or sumr_402(4) or sumr_402(5) or sumr_402(6) or sumr_402(7) or sumr_402(8) or sumr_402(9));
E(620)<=not ( sumr_403(0) or sumr_403(1) or sumr_403(2) or sumr_403(3) or sumr_403(4) or sumr_403(5) or sumr_403(6) or sumr_403(7) or sumr_403(8) or sumr_403(9));
E(619)<=not ( sumr_404(0) or sumr_404(1) or sumr_404(2) or sumr_404(3) or sumr_404(4) or sumr_404(5) or sumr_404(6) or sumr_404(7) or sumr_404(8) or sumr_404(9));
E(618)<=not ( sumr_405(0) or sumr_405(1) or sumr_405(2) or sumr_405(3) or sumr_405(4) or sumr_405(5) or sumr_405(6) or sumr_405(7) or sumr_405(8) or sumr_405(9));
E(617)<=not ( sumr_406(0) or sumr_406(1) or sumr_406(2) or sumr_406(3) or sumr_406(4) or sumr_406(5) or sumr_406(6) or sumr_406(7) or sumr_406(8) or sumr_406(9));
E(616)<=not ( sumr_407(0) or sumr_407(1) or sumr_407(2) or sumr_407(3) or sumr_407(4) or sumr_407(5) or sumr_407(6) or sumr_407(7) or sumr_407(8) or sumr_407(9));
E(615)<=not ( sumr_408(0) or sumr_408(1) or sumr_408(2) or sumr_408(3) or sumr_408(4) or sumr_408(5) or sumr_408(6) or sumr_408(7) or sumr_408(8) or sumr_408(9));
E(614)<=not ( sumr_409(0) or sumr_409(1) or sumr_409(2) or sumr_409(3) or sumr_409(4) or sumr_409(5) or sumr_409(6) or sumr_409(7) or sumr_409(8) or sumr_409(9));
E(613)<=not ( sumr_410(0) or sumr_410(1) or sumr_410(2) or sumr_410(3) or sumr_410(4) or sumr_410(5) or sumr_410(6) or sumr_410(7) or sumr_410(8) or sumr_410(9));
E(612)<=not ( sumr_411(0) or sumr_411(1) or sumr_411(2) or sumr_411(3) or sumr_411(4) or sumr_411(5) or sumr_411(6) or sumr_411(7) or sumr_411(8) or sumr_411(9));
E(611)<=not ( sumr_412(0) or sumr_412(1) or sumr_412(2) or sumr_412(3) or sumr_412(4) or sumr_412(5) or sumr_412(6) or sumr_412(7) or sumr_412(8) or sumr_412(9));
E(610)<=not ( sumr_413(0) or sumr_413(1) or sumr_413(2) or sumr_413(3) or sumr_413(4) or sumr_413(5) or sumr_413(6) or sumr_413(7) or sumr_413(8) or sumr_413(9));
E(609)<=not ( sumr_414(0) or sumr_414(1) or sumr_414(2) or sumr_414(3) or sumr_414(4) or sumr_414(5) or sumr_414(6) or sumr_414(7) or sumr_414(8) or sumr_414(9));
E(608)<=not ( sumr_415(0) or sumr_415(1) or sumr_415(2) or sumr_415(3) or sumr_415(4) or sumr_415(5) or sumr_415(6) or sumr_415(7) or sumr_415(8) or sumr_415(9));
E(607)<=not ( sumr_416(0) or sumr_416(1) or sumr_416(2) or sumr_416(3) or sumr_416(4) or sumr_416(5) or sumr_416(6) or sumr_416(7) or sumr_416(8) or sumr_416(9));
E(606)<=not ( sumr_417(0) or sumr_417(1) or sumr_417(2) or sumr_417(3) or sumr_417(4) or sumr_417(5) or sumr_417(6) or sumr_417(7) or sumr_417(8) or sumr_417(9));
E(605)<=not ( sumr_418(0) or sumr_418(1) or sumr_418(2) or sumr_418(3) or sumr_418(4) or sumr_418(5) or sumr_418(6) or sumr_418(7) or sumr_418(8) or sumr_418(9));
E(604)<=not ( sumr_419(0) or sumr_419(1) or sumr_419(2) or sumr_419(3) or sumr_419(4) or sumr_419(5) or sumr_419(6) or sumr_419(7) or sumr_419(8) or sumr_419(9));
E(603)<=not ( sumr_420(0) or sumr_420(1) or sumr_420(2) or sumr_420(3) or sumr_420(4) or sumr_420(5) or sumr_420(6) or sumr_420(7) or sumr_420(8) or sumr_420(9));
E(602)<=not ( sumr_421(0) or sumr_421(1) or sumr_421(2) or sumr_421(3) or sumr_421(4) or sumr_421(5) or sumr_421(6) or sumr_421(7) or sumr_421(8) or sumr_421(9));
E(601)<=not ( sumr_422(0) or sumr_422(1) or sumr_422(2) or sumr_422(3) or sumr_422(4) or sumr_422(5) or sumr_422(6) or sumr_422(7) or sumr_422(8) or sumr_422(9));
E(600)<=not ( sumr_423(0) or sumr_423(1) or sumr_423(2) or sumr_423(3) or sumr_423(4) or sumr_423(5) or sumr_423(6) or sumr_423(7) or sumr_423(8) or sumr_423(9));
E(599)<=not ( sumr_424(0) or sumr_424(1) or sumr_424(2) or sumr_424(3) or sumr_424(4) or sumr_424(5) or sumr_424(6) or sumr_424(7) or sumr_424(8) or sumr_424(9));
E(598)<=not ( sumr_425(0) or sumr_425(1) or sumr_425(2) or sumr_425(3) or sumr_425(4) or sumr_425(5) or sumr_425(6) or sumr_425(7) or sumr_425(8) or sumr_425(9));
E(597)<=not ( sumr_426(0) or sumr_426(1) or sumr_426(2) or sumr_426(3) or sumr_426(4) or sumr_426(5) or sumr_426(6) or sumr_426(7) or sumr_426(8) or sumr_426(9));
E(596)<=not ( sumr_427(0) or sumr_427(1) or sumr_427(2) or sumr_427(3) or sumr_427(4) or sumr_427(5) or sumr_427(6) or sumr_427(7) or sumr_427(8) or sumr_427(9));
E(595)<=not ( sumr_428(0) or sumr_428(1) or sumr_428(2) or sumr_428(3) or sumr_428(4) or sumr_428(5) or sumr_428(6) or sumr_428(7) or sumr_428(8) or sumr_428(9));
E(594)<=not ( sumr_429(0) or sumr_429(1) or sumr_429(2) or sumr_429(3) or sumr_429(4) or sumr_429(5) or sumr_429(6) or sumr_429(7) or sumr_429(8) or sumr_429(9));
E(593)<=not ( sumr_430(0) or sumr_430(1) or sumr_430(2) or sumr_430(3) or sumr_430(4) or sumr_430(5) or sumr_430(6) or sumr_430(7) or sumr_430(8) or sumr_430(9));
E(592)<=not ( sumr_431(0) or sumr_431(1) or sumr_431(2) or sumr_431(3) or sumr_431(4) or sumr_431(5) or sumr_431(6) or sumr_431(7) or sumr_431(8) or sumr_431(9));
E(591)<=not ( sumr_432(0) or sumr_432(1) or sumr_432(2) or sumr_432(3) or sumr_432(4) or sumr_432(5) or sumr_432(6) or sumr_432(7) or sumr_432(8) or sumr_432(9));
E(590)<=not ( sumr_433(0) or sumr_433(1) or sumr_433(2) or sumr_433(3) or sumr_433(4) or sumr_433(5) or sumr_433(6) or sumr_433(7) or sumr_433(8) or sumr_433(9));
E(589)<=not ( sumr_434(0) or sumr_434(1) or sumr_434(2) or sumr_434(3) or sumr_434(4) or sumr_434(5) or sumr_434(6) or sumr_434(7) or sumr_434(8) or sumr_434(9));
E(588)<=not ( sumr_435(0) or sumr_435(1) or sumr_435(2) or sumr_435(3) or sumr_435(4) or sumr_435(5) or sumr_435(6) or sumr_435(7) or sumr_435(8) or sumr_435(9));
E(587)<=not ( sumr_436(0) or sumr_436(1) or sumr_436(2) or sumr_436(3) or sumr_436(4) or sumr_436(5) or sumr_436(6) or sumr_436(7) or sumr_436(8) or sumr_436(9));
E(586)<=not ( sumr_437(0) or sumr_437(1) or sumr_437(2) or sumr_437(3) or sumr_437(4) or sumr_437(5) or sumr_437(6) or sumr_437(7) or sumr_437(8) or sumr_437(9));
E(585)<=not ( sumr_438(0) or sumr_438(1) or sumr_438(2) or sumr_438(3) or sumr_438(4) or sumr_438(5) or sumr_438(6) or sumr_438(7) or sumr_438(8) or sumr_438(9));
E(584)<=not ( sumr_439(0) or sumr_439(1) or sumr_439(2) or sumr_439(3) or sumr_439(4) or sumr_439(5) or sumr_439(6) or sumr_439(7) or sumr_439(8) or sumr_439(9));
E(583)<=not ( sumr_440(0) or sumr_440(1) or sumr_440(2) or sumr_440(3) or sumr_440(4) or sumr_440(5) or sumr_440(6) or sumr_440(7) or sumr_440(8) or sumr_440(9));
E(582)<=not ( sumr_441(0) or sumr_441(1) or sumr_441(2) or sumr_441(3) or sumr_441(4) or sumr_441(5) or sumr_441(6) or sumr_441(7) or sumr_441(8) or sumr_441(9));
E(581)<=not ( sumr_442(0) or sumr_442(1) or sumr_442(2) or sumr_442(3) or sumr_442(4) or sumr_442(5) or sumr_442(6) or sumr_442(7) or sumr_442(8) or sumr_442(9));
E(580)<=not ( sumr_443(0) or sumr_443(1) or sumr_443(2) or sumr_443(3) or sumr_443(4) or sumr_443(5) or sumr_443(6) or sumr_443(7) or sumr_443(8) or sumr_443(9));
E(579)<=not ( sumr_444(0) or sumr_444(1) or sumr_444(2) or sumr_444(3) or sumr_444(4) or sumr_444(5) or sumr_444(6) or sumr_444(7) or sumr_444(8) or sumr_444(9));
E(578)<=not ( sumr_445(0) or sumr_445(1) or sumr_445(2) or sumr_445(3) or sumr_445(4) or sumr_445(5) or sumr_445(6) or sumr_445(7) or sumr_445(8) or sumr_445(9));
E(577)<=not ( sumr_446(0) or sumr_446(1) or sumr_446(2) or sumr_446(3) or sumr_446(4) or sumr_446(5) or sumr_446(6) or sumr_446(7) or sumr_446(8) or sumr_446(9));
E(576)<=not ( sumr_447(0) or sumr_447(1) or sumr_447(2) or sumr_447(3) or sumr_447(4) or sumr_447(5) or sumr_447(6) or sumr_447(7) or sumr_447(8) or sumr_447(9));
E(575)<=not ( sumr_448(0) or sumr_448(1) or sumr_448(2) or sumr_448(3) or sumr_448(4) or sumr_448(5) or sumr_448(6) or sumr_448(7) or sumr_448(8) or sumr_448(9));
E(574)<=not ( sumr_449(0) or sumr_449(1) or sumr_449(2) or sumr_449(3) or sumr_449(4) or sumr_449(5) or sumr_449(6) or sumr_449(7) or sumr_449(8) or sumr_449(9));
E(573)<=not ( sumr_450(0) or sumr_450(1) or sumr_450(2) or sumr_450(3) or sumr_450(4) or sumr_450(5) or sumr_450(6) or sumr_450(7) or sumr_450(8) or sumr_450(9));
E(572)<=not ( sumr_451(0) or sumr_451(1) or sumr_451(2) or sumr_451(3) or sumr_451(4) or sumr_451(5) or sumr_451(6) or sumr_451(7) or sumr_451(8) or sumr_451(9));
E(571)<=not ( sumr_452(0) or sumr_452(1) or sumr_452(2) or sumr_452(3) or sumr_452(4) or sumr_452(5) or sumr_452(6) or sumr_452(7) or sumr_452(8) or sumr_452(9));
E(570)<=not ( sumr_453(0) or sumr_453(1) or sumr_453(2) or sumr_453(3) or sumr_453(4) or sumr_453(5) or sumr_453(6) or sumr_453(7) or sumr_453(8) or sumr_453(9));
E(569)<=not ( sumr_454(0) or sumr_454(1) or sumr_454(2) or sumr_454(3) or sumr_454(4) or sumr_454(5) or sumr_454(6) or sumr_454(7) or sumr_454(8) or sumr_454(9));
E(568)<=not ( sumr_455(0) or sumr_455(1) or sumr_455(2) or sumr_455(3) or sumr_455(4) or sumr_455(5) or sumr_455(6) or sumr_455(7) or sumr_455(8) or sumr_455(9));
E(567)<=not ( sumr_456(0) or sumr_456(1) or sumr_456(2) or sumr_456(3) or sumr_456(4) or sumr_456(5) or sumr_456(6) or sumr_456(7) or sumr_456(8) or sumr_456(9));
E(566)<=not ( sumr_457(0) or sumr_457(1) or sumr_457(2) or sumr_457(3) or sumr_457(4) or sumr_457(5) or sumr_457(6) or sumr_457(7) or sumr_457(8) or sumr_457(9));
E(565)<=not ( sumr_458(0) or sumr_458(1) or sumr_458(2) or sumr_458(3) or sumr_458(4) or sumr_458(5) or sumr_458(6) or sumr_458(7) or sumr_458(8) or sumr_458(9));
E(564)<=not ( sumr_459(0) or sumr_459(1) or sumr_459(2) or sumr_459(3) or sumr_459(4) or sumr_459(5) or sumr_459(6) or sumr_459(7) or sumr_459(8) or sumr_459(9));
E(563)<=not ( sumr_460(0) or sumr_460(1) or sumr_460(2) or sumr_460(3) or sumr_460(4) or sumr_460(5) or sumr_460(6) or sumr_460(7) or sumr_460(8) or sumr_460(9));
E(562)<=not ( sumr_461(0) or sumr_461(1) or sumr_461(2) or sumr_461(3) or sumr_461(4) or sumr_461(5) or sumr_461(6) or sumr_461(7) or sumr_461(8) or sumr_461(9));
E(561)<=not ( sumr_462(0) or sumr_462(1) or sumr_462(2) or sumr_462(3) or sumr_462(4) or sumr_462(5) or sumr_462(6) or sumr_462(7) or sumr_462(8) or sumr_462(9));
E(560)<=not ( sumr_463(0) or sumr_463(1) or sumr_463(2) or sumr_463(3) or sumr_463(4) or sumr_463(5) or sumr_463(6) or sumr_463(7) or sumr_463(8) or sumr_463(9));
E(559)<=not ( sumr_464(0) or sumr_464(1) or sumr_464(2) or sumr_464(3) or sumr_464(4) or sumr_464(5) or sumr_464(6) or sumr_464(7) or sumr_464(8) or sumr_464(9));
E(558)<=not ( sumr_465(0) or sumr_465(1) or sumr_465(2) or sumr_465(3) or sumr_465(4) or sumr_465(5) or sumr_465(6) or sumr_465(7) or sumr_465(8) or sumr_465(9));
E(557)<=not ( sumr_466(0) or sumr_466(1) or sumr_466(2) or sumr_466(3) or sumr_466(4) or sumr_466(5) or sumr_466(6) or sumr_466(7) or sumr_466(8) or sumr_466(9));
E(556)<=not ( sumr_467(0) or sumr_467(1) or sumr_467(2) or sumr_467(3) or sumr_467(4) or sumr_467(5) or sumr_467(6) or sumr_467(7) or sumr_467(8) or sumr_467(9));
E(555)<=not ( sumr_468(0) or sumr_468(1) or sumr_468(2) or sumr_468(3) or sumr_468(4) or sumr_468(5) or sumr_468(6) or sumr_468(7) or sumr_468(8) or sumr_468(9));
E(554)<=not ( sumr_469(0) or sumr_469(1) or sumr_469(2) or sumr_469(3) or sumr_469(4) or sumr_469(5) or sumr_469(6) or sumr_469(7) or sumr_469(8) or sumr_469(9));
E(553)<=not ( sumr_470(0) or sumr_470(1) or sumr_470(2) or sumr_470(3) or sumr_470(4) or sumr_470(5) or sumr_470(6) or sumr_470(7) or sumr_470(8) or sumr_470(9));
E(552)<=not ( sumr_471(0) or sumr_471(1) or sumr_471(2) or sumr_471(3) or sumr_471(4) or sumr_471(5) or sumr_471(6) or sumr_471(7) or sumr_471(8) or sumr_471(9));
E(551)<=not ( sumr_472(0) or sumr_472(1) or sumr_472(2) or sumr_472(3) or sumr_472(4) or sumr_472(5) or sumr_472(6) or sumr_472(7) or sumr_472(8) or sumr_472(9));
E(550)<=not ( sumr_473(0) or sumr_473(1) or sumr_473(2) or sumr_473(3) or sumr_473(4) or sumr_473(5) or sumr_473(6) or sumr_473(7) or sumr_473(8) or sumr_473(9));
E(549)<=not ( sumr_474(0) or sumr_474(1) or sumr_474(2) or sumr_474(3) or sumr_474(4) or sumr_474(5) or sumr_474(6) or sumr_474(7) or sumr_474(8) or sumr_474(9));
E(548)<=not ( sumr_475(0) or sumr_475(1) or sumr_475(2) or sumr_475(3) or sumr_475(4) or sumr_475(5) or sumr_475(6) or sumr_475(7) or sumr_475(8) or sumr_475(9));
E(547)<=not ( sumr_476(0) or sumr_476(1) or sumr_476(2) or sumr_476(3) or sumr_476(4) or sumr_476(5) or sumr_476(6) or sumr_476(7) or sumr_476(8) or sumr_476(9));
E(546)<=not ( sumr_477(0) or sumr_477(1) or sumr_477(2) or sumr_477(3) or sumr_477(4) or sumr_477(5) or sumr_477(6) or sumr_477(7) or sumr_477(8) or sumr_477(9));
E(545)<=not ( sumr_478(0) or sumr_478(1) or sumr_478(2) or sumr_478(3) or sumr_478(4) or sumr_478(5) or sumr_478(6) or sumr_478(7) or sumr_478(8) or sumr_478(9));
E(544)<=not ( sumr_479(0) or sumr_479(1) or sumr_479(2) or sumr_479(3) or sumr_479(4) or sumr_479(5) or sumr_479(6) or sumr_479(7) or sumr_479(8) or sumr_479(9));
E(543)<=not ( sumr_480(0) or sumr_480(1) or sumr_480(2) or sumr_480(3) or sumr_480(4) or sumr_480(5) or sumr_480(6) or sumr_480(7) or sumr_480(8) or sumr_480(9));
E(542)<=not ( sumr_481(0) or sumr_481(1) or sumr_481(2) or sumr_481(3) or sumr_481(4) or sumr_481(5) or sumr_481(6) or sumr_481(7) or sumr_481(8) or sumr_481(9));
E(541)<=not ( sumr_482(0) or sumr_482(1) or sumr_482(2) or sumr_482(3) or sumr_482(4) or sumr_482(5) or sumr_482(6) or sumr_482(7) or sumr_482(8) or sumr_482(9));
E(540)<=not ( sumr_483(0) or sumr_483(1) or sumr_483(2) or sumr_483(3) or sumr_483(4) or sumr_483(5) or sumr_483(6) or sumr_483(7) or sumr_483(8) or sumr_483(9));
E(539)<=not ( sumr_484(0) or sumr_484(1) or sumr_484(2) or sumr_484(3) or sumr_484(4) or sumr_484(5) or sumr_484(6) or sumr_484(7) or sumr_484(8) or sumr_484(9));
E(538)<=not ( sumr_485(0) or sumr_485(1) or sumr_485(2) or sumr_485(3) or sumr_485(4) or sumr_485(5) or sumr_485(6) or sumr_485(7) or sumr_485(8) or sumr_485(9));
E(537)<=not ( sumr_486(0) or sumr_486(1) or sumr_486(2) or sumr_486(3) or sumr_486(4) or sumr_486(5) or sumr_486(6) or sumr_486(7) or sumr_486(8) or sumr_486(9));
E(536)<=not ( sumr_487(0) or sumr_487(1) or sumr_487(2) or sumr_487(3) or sumr_487(4) or sumr_487(5) or sumr_487(6) or sumr_487(7) or sumr_487(8) or sumr_487(9));
E(535)<=not ( sumr_488(0) or sumr_488(1) or sumr_488(2) or sumr_488(3) or sumr_488(4) or sumr_488(5) or sumr_488(6) or sumr_488(7) or sumr_488(8) or sumr_488(9));
E(534)<=not ( sumr_489(0) or sumr_489(1) or sumr_489(2) or sumr_489(3) or sumr_489(4) or sumr_489(5) or sumr_489(6) or sumr_489(7) or sumr_489(8) or sumr_489(9));
E(533)<=not ( sumr_490(0) or sumr_490(1) or sumr_490(2) or sumr_490(3) or sumr_490(4) or sumr_490(5) or sumr_490(6) or sumr_490(7) or sumr_490(8) or sumr_490(9));
E(532)<=not ( sumr_491(0) or sumr_491(1) or sumr_491(2) or sumr_491(3) or sumr_491(4) or sumr_491(5) or sumr_491(6) or sumr_491(7) or sumr_491(8) or sumr_491(9));
E(531)<=not ( sumr_492(0) or sumr_492(1) or sumr_492(2) or sumr_492(3) or sumr_492(4) or sumr_492(5) or sumr_492(6) or sumr_492(7) or sumr_492(8) or sumr_492(9));
E(530)<=not ( sumr_493(0) or sumr_493(1) or sumr_493(2) or sumr_493(3) or sumr_493(4) or sumr_493(5) or sumr_493(6) or sumr_493(7) or sumr_493(8) or sumr_493(9));
E(529)<=not ( sumr_494(0) or sumr_494(1) or sumr_494(2) or sumr_494(3) or sumr_494(4) or sumr_494(5) or sumr_494(6) or sumr_494(7) or sumr_494(8) or sumr_494(9));
E(528)<=not ( sumr_495(0) or sumr_495(1) or sumr_495(2) or sumr_495(3) or sumr_495(4) or sumr_495(5) or sumr_495(6) or sumr_495(7) or sumr_495(8) or sumr_495(9));
E(527)<=not ( sumr_496(0) or sumr_496(1) or sumr_496(2) or sumr_496(3) or sumr_496(4) or sumr_496(5) or sumr_496(6) or sumr_496(7) or sumr_496(8) or sumr_496(9));
E(526)<=not ( sumr_497(0) or sumr_497(1) or sumr_497(2) or sumr_497(3) or sumr_497(4) or sumr_497(5) or sumr_497(6) or sumr_497(7) or sumr_497(8) or sumr_497(9));
E(525)<=not ( sumr_498(0) or sumr_498(1) or sumr_498(2) or sumr_498(3) or sumr_498(4) or sumr_498(5) or sumr_498(6) or sumr_498(7) or sumr_498(8) or sumr_498(9));
E(524)<=not ( sumr_499(0) or sumr_499(1) or sumr_499(2) or sumr_499(3) or sumr_499(4) or sumr_499(5) or sumr_499(6) or sumr_499(7) or sumr_499(8) or sumr_499(9));
E(523)<=not ( sumr_500(0) or sumr_500(1) or sumr_500(2) or sumr_500(3) or sumr_500(4) or sumr_500(5) or sumr_500(6) or sumr_500(7) or sumr_500(8) or sumr_500(9));
E(522)<=not ( sumr_501(0) or sumr_501(1) or sumr_501(2) or sumr_501(3) or sumr_501(4) or sumr_501(5) or sumr_501(6) or sumr_501(7) or sumr_501(8) or sumr_501(9));
E(521)<=not ( sumr_502(0) or sumr_502(1) or sumr_502(2) or sumr_502(3) or sumr_502(4) or sumr_502(5) or sumr_502(6) or sumr_502(7) or sumr_502(8) or sumr_502(9));
E(520)<=not ( sumr_503(0) or sumr_503(1) or sumr_503(2) or sumr_503(3) or sumr_503(4) or sumr_503(5) or sumr_503(6) or sumr_503(7) or sumr_503(8) or sumr_503(9));
E(519)<=not ( sumr_504(0) or sumr_504(1) or sumr_504(2) or sumr_504(3) or sumr_504(4) or sumr_504(5) or sumr_504(6) or sumr_504(7) or sumr_504(8) or sumr_504(9));
E(518)<=not ( sumr_505(0) or sumr_505(1) or sumr_505(2) or sumr_505(3) or sumr_505(4) or sumr_505(5) or sumr_505(6) or sumr_505(7) or sumr_505(8) or sumr_505(9));
E(517)<=not ( sumr_506(0) or sumr_506(1) or sumr_506(2) or sumr_506(3) or sumr_506(4) or sumr_506(5) or sumr_506(6) or sumr_506(7) or sumr_506(8) or sumr_506(9));
E(516)<=not ( sumr_507(0) or sumr_507(1) or sumr_507(2) or sumr_507(3) or sumr_507(4) or sumr_507(5) or sumr_507(6) or sumr_507(7) or sumr_507(8) or sumr_507(9));
E(515)<=not ( sumr_508(0) or sumr_508(1) or sumr_508(2) or sumr_508(3) or sumr_508(4) or sumr_508(5) or sumr_508(6) or sumr_508(7) or sumr_508(8) or sumr_508(9));
E(514)<=not ( sumr_509(0) or sumr_509(1) or sumr_509(2) or sumr_509(3) or sumr_509(4) or sumr_509(5) or sumr_509(6) or sumr_509(7) or sumr_509(8) or sumr_509(9));
E(513)<=not ( sumr_510(0) or sumr_510(1) or sumr_510(2) or sumr_510(3) or sumr_510(4) or sumr_510(5) or sumr_510(6) or sumr_510(7) or sumr_510(8) or sumr_510(9));
E(512)<=not ( sumr_511(0) or sumr_511(1) or sumr_511(2) or sumr_511(3) or sumr_511(4) or sumr_511(5) or sumr_511(6) or sumr_511(7) or sumr_511(8) or sumr_511(9));
E(511)<=not ( sumr_512(0) or sumr_512(1) or sumr_512(2) or sumr_512(3) or sumr_512(4) or sumr_512(5) or sumr_512(6) or sumr_512(7) or sumr_512(8) or sumr_512(9));
E(510)<=not ( sumr_513(0) or sumr_513(1) or sumr_513(2) or sumr_513(3) or sumr_513(4) or sumr_513(5) or sumr_513(6) or sumr_513(7) or sumr_513(8) or sumr_513(9));
E(509)<=not ( sumr_514(0) or sumr_514(1) or sumr_514(2) or sumr_514(3) or sumr_514(4) or sumr_514(5) or sumr_514(6) or sumr_514(7) or sumr_514(8) or sumr_514(9));
E(508)<=not ( sumr_515(0) or sumr_515(1) or sumr_515(2) or sumr_515(3) or sumr_515(4) or sumr_515(5) or sumr_515(6) or sumr_515(7) or sumr_515(8) or sumr_515(9));
E(507)<=not ( sumr_516(0) or sumr_516(1) or sumr_516(2) or sumr_516(3) or sumr_516(4) or sumr_516(5) or sumr_516(6) or sumr_516(7) or sumr_516(8) or sumr_516(9));
E(506)<=not ( sumr_517(0) or sumr_517(1) or sumr_517(2) or sumr_517(3) or sumr_517(4) or sumr_517(5) or sumr_517(6) or sumr_517(7) or sumr_517(8) or sumr_517(9));
E(505)<=not ( sumr_518(0) or sumr_518(1) or sumr_518(2) or sumr_518(3) or sumr_518(4) or sumr_518(5) or sumr_518(6) or sumr_518(7) or sumr_518(8) or sumr_518(9));
E(504)<=not ( sumr_519(0) or sumr_519(1) or sumr_519(2) or sumr_519(3) or sumr_519(4) or sumr_519(5) or sumr_519(6) or sumr_519(7) or sumr_519(8) or sumr_519(9));
E(503)<=not ( sumr_520(0) or sumr_520(1) or sumr_520(2) or sumr_520(3) or sumr_520(4) or sumr_520(5) or sumr_520(6) or sumr_520(7) or sumr_520(8) or sumr_520(9));
E(502)<=not ( sumr_521(0) or sumr_521(1) or sumr_521(2) or sumr_521(3) or sumr_521(4) or sumr_521(5) or sumr_521(6) or sumr_521(7) or sumr_521(8) or sumr_521(9));
E(501)<=not ( sumr_522(0) or sumr_522(1) or sumr_522(2) or sumr_522(3) or sumr_522(4) or sumr_522(5) or sumr_522(6) or sumr_522(7) or sumr_522(8) or sumr_522(9));
E(500)<=not ( sumr_523(0) or sumr_523(1) or sumr_523(2) or sumr_523(3) or sumr_523(4) or sumr_523(5) or sumr_523(6) or sumr_523(7) or sumr_523(8) or sumr_523(9));
E(499)<=not ( sumr_524(0) or sumr_524(1) or sumr_524(2) or sumr_524(3) or sumr_524(4) or sumr_524(5) or sumr_524(6) or sumr_524(7) or sumr_524(8) or sumr_524(9));
E(498)<=not ( sumr_525(0) or sumr_525(1) or sumr_525(2) or sumr_525(3) or sumr_525(4) or sumr_525(5) or sumr_525(6) or sumr_525(7) or sumr_525(8) or sumr_525(9));
E(497)<=not ( sumr_526(0) or sumr_526(1) or sumr_526(2) or sumr_526(3) or sumr_526(4) or sumr_526(5) or sumr_526(6) or sumr_526(7) or sumr_526(8) or sumr_526(9));
E(496)<=not ( sumr_527(0) or sumr_527(1) or sumr_527(2) or sumr_527(3) or sumr_527(4) or sumr_527(5) or sumr_527(6) or sumr_527(7) or sumr_527(8) or sumr_527(9));
E(495)<=not ( sumr_528(0) or sumr_528(1) or sumr_528(2) or sumr_528(3) or sumr_528(4) or sumr_528(5) or sumr_528(6) or sumr_528(7) or sumr_528(8) or sumr_528(9));
E(494)<=not ( sumr_529(0) or sumr_529(1) or sumr_529(2) or sumr_529(3) or sumr_529(4) or sumr_529(5) or sumr_529(6) or sumr_529(7) or sumr_529(8) or sumr_529(9));
E(493)<=not ( sumr_530(0) or sumr_530(1) or sumr_530(2) or sumr_530(3) or sumr_530(4) or sumr_530(5) or sumr_530(6) or sumr_530(7) or sumr_530(8) or sumr_530(9));
E(492)<=not ( sumr_531(0) or sumr_531(1) or sumr_531(2) or sumr_531(3) or sumr_531(4) or sumr_531(5) or sumr_531(6) or sumr_531(7) or sumr_531(8) or sumr_531(9));
E(491)<=not ( sumr_532(0) or sumr_532(1) or sumr_532(2) or sumr_532(3) or sumr_532(4) or sumr_532(5) or sumr_532(6) or sumr_532(7) or sumr_532(8) or sumr_532(9));
E(490)<=not ( sumr_533(0) or sumr_533(1) or sumr_533(2) or sumr_533(3) or sumr_533(4) or sumr_533(5) or sumr_533(6) or sumr_533(7) or sumr_533(8) or sumr_533(9));
E(489)<=not ( sumr_534(0) or sumr_534(1) or sumr_534(2) or sumr_534(3) or sumr_534(4) or sumr_534(5) or sumr_534(6) or sumr_534(7) or sumr_534(8) or sumr_534(9));
E(488)<=not ( sumr_535(0) or sumr_535(1) or sumr_535(2) or sumr_535(3) or sumr_535(4) or sumr_535(5) or sumr_535(6) or sumr_535(7) or sumr_535(8) or sumr_535(9));
E(487)<=not ( sumr_536(0) or sumr_536(1) or sumr_536(2) or sumr_536(3) or sumr_536(4) or sumr_536(5) or sumr_536(6) or sumr_536(7) or sumr_536(8) or sumr_536(9));
E(486)<=not ( sumr_537(0) or sumr_537(1) or sumr_537(2) or sumr_537(3) or sumr_537(4) or sumr_537(5) or sumr_537(6) or sumr_537(7) or sumr_537(8) or sumr_537(9));
E(485)<=not ( sumr_538(0) or sumr_538(1) or sumr_538(2) or sumr_538(3) or sumr_538(4) or sumr_538(5) or sumr_538(6) or sumr_538(7) or sumr_538(8) or sumr_538(9));
E(484)<=not ( sumr_539(0) or sumr_539(1) or sumr_539(2) or sumr_539(3) or sumr_539(4) or sumr_539(5) or sumr_539(6) or sumr_539(7) or sumr_539(8) or sumr_539(9));
E(483)<=not ( sumr_540(0) or sumr_540(1) or sumr_540(2) or sumr_540(3) or sumr_540(4) or sumr_540(5) or sumr_540(6) or sumr_540(7) or sumr_540(8) or sumr_540(9));
E(482)<=not ( sumr_541(0) or sumr_541(1) or sumr_541(2) or sumr_541(3) or sumr_541(4) or sumr_541(5) or sumr_541(6) or sumr_541(7) or sumr_541(8) or sumr_541(9));
E(481)<=not ( sumr_542(0) or sumr_542(1) or sumr_542(2) or sumr_542(3) or sumr_542(4) or sumr_542(5) or sumr_542(6) or sumr_542(7) or sumr_542(8) or sumr_542(9));
E(480)<=not ( sumr_543(0) or sumr_543(1) or sumr_543(2) or sumr_543(3) or sumr_543(4) or sumr_543(5) or sumr_543(6) or sumr_543(7) or sumr_543(8) or sumr_543(9));
E(479)<=not ( sumr_544(0) or sumr_544(1) or sumr_544(2) or sumr_544(3) or sumr_544(4) or sumr_544(5) or sumr_544(6) or sumr_544(7) or sumr_544(8) or sumr_544(9));
E(478)<=not ( sumr_545(0) or sumr_545(1) or sumr_545(2) or sumr_545(3) or sumr_545(4) or sumr_545(5) or sumr_545(6) or sumr_545(7) or sumr_545(8) or sumr_545(9));
E(477)<=not ( sumr_546(0) or sumr_546(1) or sumr_546(2) or sumr_546(3) or sumr_546(4) or sumr_546(5) or sumr_546(6) or sumr_546(7) or sumr_546(8) or sumr_546(9));
E(476)<=not ( sumr_547(0) or sumr_547(1) or sumr_547(2) or sumr_547(3) or sumr_547(4) or sumr_547(5) or sumr_547(6) or sumr_547(7) or sumr_547(8) or sumr_547(9));
E(475)<=not ( sumr_548(0) or sumr_548(1) or sumr_548(2) or sumr_548(3) or sumr_548(4) or sumr_548(5) or sumr_548(6) or sumr_548(7) or sumr_548(8) or sumr_548(9));
E(474)<=not ( sumr_549(0) or sumr_549(1) or sumr_549(2) or sumr_549(3) or sumr_549(4) or sumr_549(5) or sumr_549(6) or sumr_549(7) or sumr_549(8) or sumr_549(9));
E(473)<=not ( sumr_550(0) or sumr_550(1) or sumr_550(2) or sumr_550(3) or sumr_550(4) or sumr_550(5) or sumr_550(6) or sumr_550(7) or sumr_550(8) or sumr_550(9));
E(472)<=not ( sumr_551(0) or sumr_551(1) or sumr_551(2) or sumr_551(3) or sumr_551(4) or sumr_551(5) or sumr_551(6) or sumr_551(7) or sumr_551(8) or sumr_551(9));
E(471)<=not ( sumr_552(0) or sumr_552(1) or sumr_552(2) or sumr_552(3) or sumr_552(4) or sumr_552(5) or sumr_552(6) or sumr_552(7) or sumr_552(8) or sumr_552(9));
E(470)<=not ( sumr_553(0) or sumr_553(1) or sumr_553(2) or sumr_553(3) or sumr_553(4) or sumr_553(5) or sumr_553(6) or sumr_553(7) or sumr_553(8) or sumr_553(9));
E(469)<=not ( sumr_554(0) or sumr_554(1) or sumr_554(2) or sumr_554(3) or sumr_554(4) or sumr_554(5) or sumr_554(6) or sumr_554(7) or sumr_554(8) or sumr_554(9));
E(468)<=not ( sumr_555(0) or sumr_555(1) or sumr_555(2) or sumr_555(3) or sumr_555(4) or sumr_555(5) or sumr_555(6) or sumr_555(7) or sumr_555(8) or sumr_555(9));
E(467)<=not ( sumr_556(0) or sumr_556(1) or sumr_556(2) or sumr_556(3) or sumr_556(4) or sumr_556(5) or sumr_556(6) or sumr_556(7) or sumr_556(8) or sumr_556(9));
E(466)<=not ( sumr_557(0) or sumr_557(1) or sumr_557(2) or sumr_557(3) or sumr_557(4) or sumr_557(5) or sumr_557(6) or sumr_557(7) or sumr_557(8) or sumr_557(9));
E(465)<=not ( sumr_558(0) or sumr_558(1) or sumr_558(2) or sumr_558(3) or sumr_558(4) or sumr_558(5) or sumr_558(6) or sumr_558(7) or sumr_558(8) or sumr_558(9));
E(464)<=not ( sumr_559(0) or sumr_559(1) or sumr_559(2) or sumr_559(3) or sumr_559(4) or sumr_559(5) or sumr_559(6) or sumr_559(7) or sumr_559(8) or sumr_559(9));
E(463)<=not ( sumr_560(0) or sumr_560(1) or sumr_560(2) or sumr_560(3) or sumr_560(4) or sumr_560(5) or sumr_560(6) or sumr_560(7) or sumr_560(8) or sumr_560(9));
E(462)<=not ( sumr_561(0) or sumr_561(1) or sumr_561(2) or sumr_561(3) or sumr_561(4) or sumr_561(5) or sumr_561(6) or sumr_561(7) or sumr_561(8) or sumr_561(9));
E(461)<=not ( sumr_562(0) or sumr_562(1) or sumr_562(2) or sumr_562(3) or sumr_562(4) or sumr_562(5) or sumr_562(6) or sumr_562(7) or sumr_562(8) or sumr_562(9));
E(460)<=not ( sumr_563(0) or sumr_563(1) or sumr_563(2) or sumr_563(3) or sumr_563(4) or sumr_563(5) or sumr_563(6) or sumr_563(7) or sumr_563(8) or sumr_563(9));
E(459)<=not ( sumr_564(0) or sumr_564(1) or sumr_564(2) or sumr_564(3) or sumr_564(4) or sumr_564(5) or sumr_564(6) or sumr_564(7) or sumr_564(8) or sumr_564(9));
E(458)<=not ( sumr_565(0) or sumr_565(1) or sumr_565(2) or sumr_565(3) or sumr_565(4) or sumr_565(5) or sumr_565(6) or sumr_565(7) or sumr_565(8) or sumr_565(9));
E(457)<=not ( sumr_566(0) or sumr_566(1) or sumr_566(2) or sumr_566(3) or sumr_566(4) or sumr_566(5) or sumr_566(6) or sumr_566(7) or sumr_566(8) or sumr_566(9));
E(456)<=not ( sumr_567(0) or sumr_567(1) or sumr_567(2) or sumr_567(3) or sumr_567(4) or sumr_567(5) or sumr_567(6) or sumr_567(7) or sumr_567(8) or sumr_567(9));
E(455)<=not ( sumr_568(0) or sumr_568(1) or sumr_568(2) or sumr_568(3) or sumr_568(4) or sumr_568(5) or sumr_568(6) or sumr_568(7) or sumr_568(8) or sumr_568(9));
E(454)<=not ( sumr_569(0) or sumr_569(1) or sumr_569(2) or sumr_569(3) or sumr_569(4) or sumr_569(5) or sumr_569(6) or sumr_569(7) or sumr_569(8) or sumr_569(9));
E(453)<=not ( sumr_570(0) or sumr_570(1) or sumr_570(2) or sumr_570(3) or sumr_570(4) or sumr_570(5) or sumr_570(6) or sumr_570(7) or sumr_570(8) or sumr_570(9));
E(452)<=not ( sumr_571(0) or sumr_571(1) or sumr_571(2) or sumr_571(3) or sumr_571(4) or sumr_571(5) or sumr_571(6) or sumr_571(7) or sumr_571(8) or sumr_571(9));
E(451)<=not ( sumr_572(0) or sumr_572(1) or sumr_572(2) or sumr_572(3) or sumr_572(4) or sumr_572(5) or sumr_572(6) or sumr_572(7) or sumr_572(8) or sumr_572(9));
E(450)<=not ( sumr_573(0) or sumr_573(1) or sumr_573(2) or sumr_573(3) or sumr_573(4) or sumr_573(5) or sumr_573(6) or sumr_573(7) or sumr_573(8) or sumr_573(9));
E(449)<=not ( sumr_574(0) or sumr_574(1) or sumr_574(2) or sumr_574(3) or sumr_574(4) or sumr_574(5) or sumr_574(6) or sumr_574(7) or sumr_574(8) or sumr_574(9));
E(448)<=not ( sumr_575(0) or sumr_575(1) or sumr_575(2) or sumr_575(3) or sumr_575(4) or sumr_575(5) or sumr_575(6) or sumr_575(7) or sumr_575(8) or sumr_575(9));
E(447)<=not ( sumr_576(0) or sumr_576(1) or sumr_576(2) or sumr_576(3) or sumr_576(4) or sumr_576(5) or sumr_576(6) or sumr_576(7) or sumr_576(8) or sumr_576(9));
E(446)<=not ( sumr_577(0) or sumr_577(1) or sumr_577(2) or sumr_577(3) or sumr_577(4) or sumr_577(5) or sumr_577(6) or sumr_577(7) or sumr_577(8) or sumr_577(9));
E(445)<=not ( sumr_578(0) or sumr_578(1) or sumr_578(2) or sumr_578(3) or sumr_578(4) or sumr_578(5) or sumr_578(6) or sumr_578(7) or sumr_578(8) or sumr_578(9));
E(444)<=not ( sumr_579(0) or sumr_579(1) or sumr_579(2) or sumr_579(3) or sumr_579(4) or sumr_579(5) or sumr_579(6) or sumr_579(7) or sumr_579(8) or sumr_579(9));
E(443)<=not ( sumr_580(0) or sumr_580(1) or sumr_580(2) or sumr_580(3) or sumr_580(4) or sumr_580(5) or sumr_580(6) or sumr_580(7) or sumr_580(8) or sumr_580(9));
E(442)<=not ( sumr_581(0) or sumr_581(1) or sumr_581(2) or sumr_581(3) or sumr_581(4) or sumr_581(5) or sumr_581(6) or sumr_581(7) or sumr_581(8) or sumr_581(9));
E(441)<=not ( sumr_582(0) or sumr_582(1) or sumr_582(2) or sumr_582(3) or sumr_582(4) or sumr_582(5) or sumr_582(6) or sumr_582(7) or sumr_582(8) or sumr_582(9));
E(440)<=not ( sumr_583(0) or sumr_583(1) or sumr_583(2) or sumr_583(3) or sumr_583(4) or sumr_583(5) or sumr_583(6) or sumr_583(7) or sumr_583(8) or sumr_583(9));
E(439)<=not ( sumr_584(0) or sumr_584(1) or sumr_584(2) or sumr_584(3) or sumr_584(4) or sumr_584(5) or sumr_584(6) or sumr_584(7) or sumr_584(8) or sumr_584(9));
E(438)<=not ( sumr_585(0) or sumr_585(1) or sumr_585(2) or sumr_585(3) or sumr_585(4) or sumr_585(5) or sumr_585(6) or sumr_585(7) or sumr_585(8) or sumr_585(9));
E(437)<=not ( sumr_586(0) or sumr_586(1) or sumr_586(2) or sumr_586(3) or sumr_586(4) or sumr_586(5) or sumr_586(6) or sumr_586(7) or sumr_586(8) or sumr_586(9));
E(436)<=not ( sumr_587(0) or sumr_587(1) or sumr_587(2) or sumr_587(3) or sumr_587(4) or sumr_587(5) or sumr_587(6) or sumr_587(7) or sumr_587(8) or sumr_587(9));
E(435)<=not ( sumr_588(0) or sumr_588(1) or sumr_588(2) or sumr_588(3) or sumr_588(4) or sumr_588(5) or sumr_588(6) or sumr_588(7) or sumr_588(8) or sumr_588(9));
E(434)<=not ( sumr_589(0) or sumr_589(1) or sumr_589(2) or sumr_589(3) or sumr_589(4) or sumr_589(5) or sumr_589(6) or sumr_589(7) or sumr_589(8) or sumr_589(9));
E(433)<=not ( sumr_590(0) or sumr_590(1) or sumr_590(2) or sumr_590(3) or sumr_590(4) or sumr_590(5) or sumr_590(6) or sumr_590(7) or sumr_590(8) or sumr_590(9));
E(432)<=not ( sumr_591(0) or sumr_591(1) or sumr_591(2) or sumr_591(3) or sumr_591(4) or sumr_591(5) or sumr_591(6) or sumr_591(7) or sumr_591(8) or sumr_591(9));
E(431)<=not ( sumr_592(0) or sumr_592(1) or sumr_592(2) or sumr_592(3) or sumr_592(4) or sumr_592(5) or sumr_592(6) or sumr_592(7) or sumr_592(8) or sumr_592(9));
E(430)<=not ( sumr_593(0) or sumr_593(1) or sumr_593(2) or sumr_593(3) or sumr_593(4) or sumr_593(5) or sumr_593(6) or sumr_593(7) or sumr_593(8) or sumr_593(9));
E(429)<=not ( sumr_594(0) or sumr_594(1) or sumr_594(2) or sumr_594(3) or sumr_594(4) or sumr_594(5) or sumr_594(6) or sumr_594(7) or sumr_594(8) or sumr_594(9));
E(428)<=not ( sumr_595(0) or sumr_595(1) or sumr_595(2) or sumr_595(3) or sumr_595(4) or sumr_595(5) or sumr_595(6) or sumr_595(7) or sumr_595(8) or sumr_595(9));
E(427)<=not ( sumr_596(0) or sumr_596(1) or sumr_596(2) or sumr_596(3) or sumr_596(4) or sumr_596(5) or sumr_596(6) or sumr_596(7) or sumr_596(8) or sumr_596(9));
E(426)<=not ( sumr_597(0) or sumr_597(1) or sumr_597(2) or sumr_597(3) or sumr_597(4) or sumr_597(5) or sumr_597(6) or sumr_597(7) or sumr_597(8) or sumr_597(9));
E(425)<=not ( sumr_598(0) or sumr_598(1) or sumr_598(2) or sumr_598(3) or sumr_598(4) or sumr_598(5) or sumr_598(6) or sumr_598(7) or sumr_598(8) or sumr_598(9));
E(424)<=not ( sumr_599(0) or sumr_599(1) or sumr_599(2) or sumr_599(3) or sumr_599(4) or sumr_599(5) or sumr_599(6) or sumr_599(7) or sumr_599(8) or sumr_599(9));
E(423)<=not ( sumr_600(0) or sumr_600(1) or sumr_600(2) or sumr_600(3) or sumr_600(4) or sumr_600(5) or sumr_600(6) or sumr_600(7) or sumr_600(8) or sumr_600(9));
E(422)<=not ( sumr_601(0) or sumr_601(1) or sumr_601(2) or sumr_601(3) or sumr_601(4) or sumr_601(5) or sumr_601(6) or sumr_601(7) or sumr_601(8) or sumr_601(9));
E(421)<=not ( sumr_602(0) or sumr_602(1) or sumr_602(2) or sumr_602(3) or sumr_602(4) or sumr_602(5) or sumr_602(6) or sumr_602(7) or sumr_602(8) or sumr_602(9));
E(420)<=not ( sumr_603(0) or sumr_603(1) or sumr_603(2) or sumr_603(3) or sumr_603(4) or sumr_603(5) or sumr_603(6) or sumr_603(7) or sumr_603(8) or sumr_603(9));
E(419)<=not ( sumr_604(0) or sumr_604(1) or sumr_604(2) or sumr_604(3) or sumr_604(4) or sumr_604(5) or sumr_604(6) or sumr_604(7) or sumr_604(8) or sumr_604(9));
E(418)<=not ( sumr_605(0) or sumr_605(1) or sumr_605(2) or sumr_605(3) or sumr_605(4) or sumr_605(5) or sumr_605(6) or sumr_605(7) or sumr_605(8) or sumr_605(9));
E(417)<=not ( sumr_606(0) or sumr_606(1) or sumr_606(2) or sumr_606(3) or sumr_606(4) or sumr_606(5) or sumr_606(6) or sumr_606(7) or sumr_606(8) or sumr_606(9));
E(416)<=not ( sumr_607(0) or sumr_607(1) or sumr_607(2) or sumr_607(3) or sumr_607(4) or sumr_607(5) or sumr_607(6) or sumr_607(7) or sumr_607(8) or sumr_607(9));
E(415)<=not ( sumr_608(0) or sumr_608(1) or sumr_608(2) or sumr_608(3) or sumr_608(4) or sumr_608(5) or sumr_608(6) or sumr_608(7) or sumr_608(8) or sumr_608(9));
E(414)<=not ( sumr_609(0) or sumr_609(1) or sumr_609(2) or sumr_609(3) or sumr_609(4) or sumr_609(5) or sumr_609(6) or sumr_609(7) or sumr_609(8) or sumr_609(9));
E(413)<=not ( sumr_610(0) or sumr_610(1) or sumr_610(2) or sumr_610(3) or sumr_610(4) or sumr_610(5) or sumr_610(6) or sumr_610(7) or sumr_610(8) or sumr_610(9));
E(412)<=not ( sumr_611(0) or sumr_611(1) or sumr_611(2) or sumr_611(3) or sumr_611(4) or sumr_611(5) or sumr_611(6) or sumr_611(7) or sumr_611(8) or sumr_611(9));
E(411)<=not ( sumr_612(0) or sumr_612(1) or sumr_612(2) or sumr_612(3) or sumr_612(4) or sumr_612(5) or sumr_612(6) or sumr_612(7) or sumr_612(8) or sumr_612(9));
E(410)<=not ( sumr_613(0) or sumr_613(1) or sumr_613(2) or sumr_613(3) or sumr_613(4) or sumr_613(5) or sumr_613(6) or sumr_613(7) or sumr_613(8) or sumr_613(9));
E(409)<=not ( sumr_614(0) or sumr_614(1) or sumr_614(2) or sumr_614(3) or sumr_614(4) or sumr_614(5) or sumr_614(6) or sumr_614(7) or sumr_614(8) or sumr_614(9));
E(408)<=not ( sumr_615(0) or sumr_615(1) or sumr_615(2) or sumr_615(3) or sumr_615(4) or sumr_615(5) or sumr_615(6) or sumr_615(7) or sumr_615(8) or sumr_615(9));
E(407)<=not ( sumr_616(0) or sumr_616(1) or sumr_616(2) or sumr_616(3) or sumr_616(4) or sumr_616(5) or sumr_616(6) or sumr_616(7) or sumr_616(8) or sumr_616(9));
E(406)<=not ( sumr_617(0) or sumr_617(1) or sumr_617(2) or sumr_617(3) or sumr_617(4) or sumr_617(5) or sumr_617(6) or sumr_617(7) or sumr_617(8) or sumr_617(9));
E(405)<=not ( sumr_618(0) or sumr_618(1) or sumr_618(2) or sumr_618(3) or sumr_618(4) or sumr_618(5) or sumr_618(6) or sumr_618(7) or sumr_618(8) or sumr_618(9));
E(404)<=not ( sumr_619(0) or sumr_619(1) or sumr_619(2) or sumr_619(3) or sumr_619(4) or sumr_619(5) or sumr_619(6) or sumr_619(7) or sumr_619(8) or sumr_619(9));
E(403)<=not ( sumr_620(0) or sumr_620(1) or sumr_620(2) or sumr_620(3) or sumr_620(4) or sumr_620(5) or sumr_620(6) or sumr_620(7) or sumr_620(8) or sumr_620(9));
E(402)<=not ( sumr_621(0) or sumr_621(1) or sumr_621(2) or sumr_621(3) or sumr_621(4) or sumr_621(5) or sumr_621(6) or sumr_621(7) or sumr_621(8) or sumr_621(9));
E(401)<=not ( sumr_622(0) or sumr_622(1) or sumr_622(2) or sumr_622(3) or sumr_622(4) or sumr_622(5) or sumr_622(6) or sumr_622(7) or sumr_622(8) or sumr_622(9));
E(400)<=not ( sumr_623(0) or sumr_623(1) or sumr_623(2) or sumr_623(3) or sumr_623(4) or sumr_623(5) or sumr_623(6) or sumr_623(7) or sumr_623(8) or sumr_623(9));
E(399)<=not ( sumr_624(0) or sumr_624(1) or sumr_624(2) or sumr_624(3) or sumr_624(4) or sumr_624(5) or sumr_624(6) or sumr_624(7) or sumr_624(8) or sumr_624(9));
E(398)<=not ( sumr_625(0) or sumr_625(1) or sumr_625(2) or sumr_625(3) or sumr_625(4) or sumr_625(5) or sumr_625(6) or sumr_625(7) or sumr_625(8) or sumr_625(9));
E(397)<=not ( sumr_626(0) or sumr_626(1) or sumr_626(2) or sumr_626(3) or sumr_626(4) or sumr_626(5) or sumr_626(6) or sumr_626(7) or sumr_626(8) or sumr_626(9));
E(396)<=not ( sumr_627(0) or sumr_627(1) or sumr_627(2) or sumr_627(3) or sumr_627(4) or sumr_627(5) or sumr_627(6) or sumr_627(7) or sumr_627(8) or sumr_627(9));
E(395)<=not ( sumr_628(0) or sumr_628(1) or sumr_628(2) or sumr_628(3) or sumr_628(4) or sumr_628(5) or sumr_628(6) or sumr_628(7) or sumr_628(8) or sumr_628(9));
E(394)<=not ( sumr_629(0) or sumr_629(1) or sumr_629(2) or sumr_629(3) or sumr_629(4) or sumr_629(5) or sumr_629(6) or sumr_629(7) or sumr_629(8) or sumr_629(9));
E(393)<=not ( sumr_630(0) or sumr_630(1) or sumr_630(2) or sumr_630(3) or sumr_630(4) or sumr_630(5) or sumr_630(6) or sumr_630(7) or sumr_630(8) or sumr_630(9));
E(392)<=not ( sumr_631(0) or sumr_631(1) or sumr_631(2) or sumr_631(3) or sumr_631(4) or sumr_631(5) or sumr_631(6) or sumr_631(7) or sumr_631(8) or sumr_631(9));
E(391)<=not ( sumr_632(0) or sumr_632(1) or sumr_632(2) or sumr_632(3) or sumr_632(4) or sumr_632(5) or sumr_632(6) or sumr_632(7) or sumr_632(8) or sumr_632(9));
E(390)<=not ( sumr_633(0) or sumr_633(1) or sumr_633(2) or sumr_633(3) or sumr_633(4) or sumr_633(5) or sumr_633(6) or sumr_633(7) or sumr_633(8) or sumr_633(9));
E(389)<=not ( sumr_634(0) or sumr_634(1) or sumr_634(2) or sumr_634(3) or sumr_634(4) or sumr_634(5) or sumr_634(6) or sumr_634(7) or sumr_634(8) or sumr_634(9));
E(388)<=not ( sumr_635(0) or sumr_635(1) or sumr_635(2) or sumr_635(3) or sumr_635(4) or sumr_635(5) or sumr_635(6) or sumr_635(7) or sumr_635(8) or sumr_635(9));
E(387)<=not ( sumr_636(0) or sumr_636(1) or sumr_636(2) or sumr_636(3) or sumr_636(4) or sumr_636(5) or sumr_636(6) or sumr_636(7) or sumr_636(8) or sumr_636(9));
E(386)<=not ( sumr_637(0) or sumr_637(1) or sumr_637(2) or sumr_637(3) or sumr_637(4) or sumr_637(5) or sumr_637(6) or sumr_637(7) or sumr_637(8) or sumr_637(9));
E(385)<=not ( sumr_638(0) or sumr_638(1) or sumr_638(2) or sumr_638(3) or sumr_638(4) or sumr_638(5) or sumr_638(6) or sumr_638(7) or sumr_638(8) or sumr_638(9));
E(384)<=not ( sumr_639(0) or sumr_639(1) or sumr_639(2) or sumr_639(3) or sumr_639(4) or sumr_639(5) or sumr_639(6) or sumr_639(7) or sumr_639(8) or sumr_639(9));
E(383)<=not ( sumr_640(0) or sumr_640(1) or sumr_640(2) or sumr_640(3) or sumr_640(4) or sumr_640(5) or sumr_640(6) or sumr_640(7) or sumr_640(8) or sumr_640(9));
E(382)<=not ( sumr_641(0) or sumr_641(1) or sumr_641(2) or sumr_641(3) or sumr_641(4) or sumr_641(5) or sumr_641(6) or sumr_641(7) or sumr_641(8) or sumr_641(9));
E(381)<=not ( sumr_642(0) or sumr_642(1) or sumr_642(2) or sumr_642(3) or sumr_642(4) or sumr_642(5) or sumr_642(6) or sumr_642(7) or sumr_642(8) or sumr_642(9));
E(380)<=not ( sumr_643(0) or sumr_643(1) or sumr_643(2) or sumr_643(3) or sumr_643(4) or sumr_643(5) or sumr_643(6) or sumr_643(7) or sumr_643(8) or sumr_643(9));
E(379)<=not ( sumr_644(0) or sumr_644(1) or sumr_644(2) or sumr_644(3) or sumr_644(4) or sumr_644(5) or sumr_644(6) or sumr_644(7) or sumr_644(8) or sumr_644(9));
E(378)<=not ( sumr_645(0) or sumr_645(1) or sumr_645(2) or sumr_645(3) or sumr_645(4) or sumr_645(5) or sumr_645(6) or sumr_645(7) or sumr_645(8) or sumr_645(9));
E(377)<=not ( sumr_646(0) or sumr_646(1) or sumr_646(2) or sumr_646(3) or sumr_646(4) or sumr_646(5) or sumr_646(6) or sumr_646(7) or sumr_646(8) or sumr_646(9));
E(376)<=not ( sumr_647(0) or sumr_647(1) or sumr_647(2) or sumr_647(3) or sumr_647(4) or sumr_647(5) or sumr_647(6) or sumr_647(7) or sumr_647(8) or sumr_647(9));
E(375)<=not ( sumr_648(0) or sumr_648(1) or sumr_648(2) or sumr_648(3) or sumr_648(4) or sumr_648(5) or sumr_648(6) or sumr_648(7) or sumr_648(8) or sumr_648(9));
E(374)<=not ( sumr_649(0) or sumr_649(1) or sumr_649(2) or sumr_649(3) or sumr_649(4) or sumr_649(5) or sumr_649(6) or sumr_649(7) or sumr_649(8) or sumr_649(9));
E(373)<=not ( sumr_650(0) or sumr_650(1) or sumr_650(2) or sumr_650(3) or sumr_650(4) or sumr_650(5) or sumr_650(6) or sumr_650(7) or sumr_650(8) or sumr_650(9));
E(372)<=not ( sumr_651(0) or sumr_651(1) or sumr_651(2) or sumr_651(3) or sumr_651(4) or sumr_651(5) or sumr_651(6) or sumr_651(7) or sumr_651(8) or sumr_651(9));
E(371)<=not ( sumr_652(0) or sumr_652(1) or sumr_652(2) or sumr_652(3) or sumr_652(4) or sumr_652(5) or sumr_652(6) or sumr_652(7) or sumr_652(8) or sumr_652(9));
E(370)<=not ( sumr_653(0) or sumr_653(1) or sumr_653(2) or sumr_653(3) or sumr_653(4) or sumr_653(5) or sumr_653(6) or sumr_653(7) or sumr_653(8) or sumr_653(9));
E(369)<=not ( sumr_654(0) or sumr_654(1) or sumr_654(2) or sumr_654(3) or sumr_654(4) or sumr_654(5) or sumr_654(6) or sumr_654(7) or sumr_654(8) or sumr_654(9));
E(368)<=not ( sumr_655(0) or sumr_655(1) or sumr_655(2) or sumr_655(3) or sumr_655(4) or sumr_655(5) or sumr_655(6) or sumr_655(7) or sumr_655(8) or sumr_655(9));
E(367)<=not ( sumr_656(0) or sumr_656(1) or sumr_656(2) or sumr_656(3) or sumr_656(4) or sumr_656(5) or sumr_656(6) or sumr_656(7) or sumr_656(8) or sumr_656(9));
E(366)<=not ( sumr_657(0) or sumr_657(1) or sumr_657(2) or sumr_657(3) or sumr_657(4) or sumr_657(5) or sumr_657(6) or sumr_657(7) or sumr_657(8) or sumr_657(9));
E(365)<=not ( sumr_658(0) or sumr_658(1) or sumr_658(2) or sumr_658(3) or sumr_658(4) or sumr_658(5) or sumr_658(6) or sumr_658(7) or sumr_658(8) or sumr_658(9));
E(364)<=not ( sumr_659(0) or sumr_659(1) or sumr_659(2) or sumr_659(3) or sumr_659(4) or sumr_659(5) or sumr_659(6) or sumr_659(7) or sumr_659(8) or sumr_659(9));
E(363)<=not ( sumr_660(0) or sumr_660(1) or sumr_660(2) or sumr_660(3) or sumr_660(4) or sumr_660(5) or sumr_660(6) or sumr_660(7) or sumr_660(8) or sumr_660(9));
E(362)<=not ( sumr_661(0) or sumr_661(1) or sumr_661(2) or sumr_661(3) or sumr_661(4) or sumr_661(5) or sumr_661(6) or sumr_661(7) or sumr_661(8) or sumr_661(9));
E(361)<=not ( sumr_662(0) or sumr_662(1) or sumr_662(2) or sumr_662(3) or sumr_662(4) or sumr_662(5) or sumr_662(6) or sumr_662(7) or sumr_662(8) or sumr_662(9));
E(360)<=not ( sumr_663(0) or sumr_663(1) or sumr_663(2) or sumr_663(3) or sumr_663(4) or sumr_663(5) or sumr_663(6) or sumr_663(7) or sumr_663(8) or sumr_663(9));
E(359)<=not ( sumr_664(0) or sumr_664(1) or sumr_664(2) or sumr_664(3) or sumr_664(4) or sumr_664(5) or sumr_664(6) or sumr_664(7) or sumr_664(8) or sumr_664(9));
E(358)<=not ( sumr_665(0) or sumr_665(1) or sumr_665(2) or sumr_665(3) or sumr_665(4) or sumr_665(5) or sumr_665(6) or sumr_665(7) or sumr_665(8) or sumr_665(9));
E(357)<=not ( sumr_666(0) or sumr_666(1) or sumr_666(2) or sumr_666(3) or sumr_666(4) or sumr_666(5) or sumr_666(6) or sumr_666(7) or sumr_666(8) or sumr_666(9));
E(356)<=not ( sumr_667(0) or sumr_667(1) or sumr_667(2) or sumr_667(3) or sumr_667(4) or sumr_667(5) or sumr_667(6) or sumr_667(7) or sumr_667(8) or sumr_667(9));
E(355)<=not ( sumr_668(0) or sumr_668(1) or sumr_668(2) or sumr_668(3) or sumr_668(4) or sumr_668(5) or sumr_668(6) or sumr_668(7) or sumr_668(8) or sumr_668(9));
E(354)<=not ( sumr_669(0) or sumr_669(1) or sumr_669(2) or sumr_669(3) or sumr_669(4) or sumr_669(5) or sumr_669(6) or sumr_669(7) or sumr_669(8) or sumr_669(9));
E(353)<=not ( sumr_670(0) or sumr_670(1) or sumr_670(2) or sumr_670(3) or sumr_670(4) or sumr_670(5) or sumr_670(6) or sumr_670(7) or sumr_670(8) or sumr_670(9));
E(352)<=not ( sumr_671(0) or sumr_671(1) or sumr_671(2) or sumr_671(3) or sumr_671(4) or sumr_671(5) or sumr_671(6) or sumr_671(7) or sumr_671(8) or sumr_671(9));
E(351)<=not ( sumr_672(0) or sumr_672(1) or sumr_672(2) or sumr_672(3) or sumr_672(4) or sumr_672(5) or sumr_672(6) or sumr_672(7) or sumr_672(8) or sumr_672(9));
E(350)<=not ( sumr_673(0) or sumr_673(1) or sumr_673(2) or sumr_673(3) or sumr_673(4) or sumr_673(5) or sumr_673(6) or sumr_673(7) or sumr_673(8) or sumr_673(9));
E(349)<=not ( sumr_674(0) or sumr_674(1) or sumr_674(2) or sumr_674(3) or sumr_674(4) or sumr_674(5) or sumr_674(6) or sumr_674(7) or sumr_674(8) or sumr_674(9));
E(348)<=not ( sumr_675(0) or sumr_675(1) or sumr_675(2) or sumr_675(3) or sumr_675(4) or sumr_675(5) or sumr_675(6) or sumr_675(7) or sumr_675(8) or sumr_675(9));
E(347)<=not ( sumr_676(0) or sumr_676(1) or sumr_676(2) or sumr_676(3) or sumr_676(4) or sumr_676(5) or sumr_676(6) or sumr_676(7) or sumr_676(8) or sumr_676(9));
E(346)<=not ( sumr_677(0) or sumr_677(1) or sumr_677(2) or sumr_677(3) or sumr_677(4) or sumr_677(5) or sumr_677(6) or sumr_677(7) or sumr_677(8) or sumr_677(9));
E(345)<=not ( sumr_678(0) or sumr_678(1) or sumr_678(2) or sumr_678(3) or sumr_678(4) or sumr_678(5) or sumr_678(6) or sumr_678(7) or sumr_678(8) or sumr_678(9));
E(344)<=not ( sumr_679(0) or sumr_679(1) or sumr_679(2) or sumr_679(3) or sumr_679(4) or sumr_679(5) or sumr_679(6) or sumr_679(7) or sumr_679(8) or sumr_679(9));
E(343)<=not ( sumr_680(0) or sumr_680(1) or sumr_680(2) or sumr_680(3) or sumr_680(4) or sumr_680(5) or sumr_680(6) or sumr_680(7) or sumr_680(8) or sumr_680(9));
E(342)<=not ( sumr_681(0) or sumr_681(1) or sumr_681(2) or sumr_681(3) or sumr_681(4) or sumr_681(5) or sumr_681(6) or sumr_681(7) or sumr_681(8) or sumr_681(9));
E(341)<=not ( sumr_682(0) or sumr_682(1) or sumr_682(2) or sumr_682(3) or sumr_682(4) or sumr_682(5) or sumr_682(6) or sumr_682(7) or sumr_682(8) or sumr_682(9));
E(340)<=not ( sumr_683(0) or sumr_683(1) or sumr_683(2) or sumr_683(3) or sumr_683(4) or sumr_683(5) or sumr_683(6) or sumr_683(7) or sumr_683(8) or sumr_683(9));
E(339)<=not ( sumr_684(0) or sumr_684(1) or sumr_684(2) or sumr_684(3) or sumr_684(4) or sumr_684(5) or sumr_684(6) or sumr_684(7) or sumr_684(8) or sumr_684(9));
E(338)<=not ( sumr_685(0) or sumr_685(1) or sumr_685(2) or sumr_685(3) or sumr_685(4) or sumr_685(5) or sumr_685(6) or sumr_685(7) or sumr_685(8) or sumr_685(9));
E(337)<=not ( sumr_686(0) or sumr_686(1) or sumr_686(2) or sumr_686(3) or sumr_686(4) or sumr_686(5) or sumr_686(6) or sumr_686(7) or sumr_686(8) or sumr_686(9));
E(336)<=not ( sumr_687(0) or sumr_687(1) or sumr_687(2) or sumr_687(3) or sumr_687(4) or sumr_687(5) or sumr_687(6) or sumr_687(7) or sumr_687(8) or sumr_687(9));
E(335)<=not ( sumr_688(0) or sumr_688(1) or sumr_688(2) or sumr_688(3) or sumr_688(4) or sumr_688(5) or sumr_688(6) or sumr_688(7) or sumr_688(8) or sumr_688(9));
E(334)<=not ( sumr_689(0) or sumr_689(1) or sumr_689(2) or sumr_689(3) or sumr_689(4) or sumr_689(5) or sumr_689(6) or sumr_689(7) or sumr_689(8) or sumr_689(9));
E(333)<=not ( sumr_690(0) or sumr_690(1) or sumr_690(2) or sumr_690(3) or sumr_690(4) or sumr_690(5) or sumr_690(6) or sumr_690(7) or sumr_690(8) or sumr_690(9));
E(332)<=not ( sumr_691(0) or sumr_691(1) or sumr_691(2) or sumr_691(3) or sumr_691(4) or sumr_691(5) or sumr_691(6) or sumr_691(7) or sumr_691(8) or sumr_691(9));
E(331)<=not ( sumr_692(0) or sumr_692(1) or sumr_692(2) or sumr_692(3) or sumr_692(4) or sumr_692(5) or sumr_692(6) or sumr_692(7) or sumr_692(8) or sumr_692(9));
E(330)<=not ( sumr_693(0) or sumr_693(1) or sumr_693(2) or sumr_693(3) or sumr_693(4) or sumr_693(5) or sumr_693(6) or sumr_693(7) or sumr_693(8) or sumr_693(9));
E(329)<=not ( sumr_694(0) or sumr_694(1) or sumr_694(2) or sumr_694(3) or sumr_694(4) or sumr_694(5) or sumr_694(6) or sumr_694(7) or sumr_694(8) or sumr_694(9));
E(328)<=not ( sumr_695(0) or sumr_695(1) or sumr_695(2) or sumr_695(3) or sumr_695(4) or sumr_695(5) or sumr_695(6) or sumr_695(7) or sumr_695(8) or sumr_695(9));
E(327)<=not ( sumr_696(0) or sumr_696(1) or sumr_696(2) or sumr_696(3) or sumr_696(4) or sumr_696(5) or sumr_696(6) or sumr_696(7) or sumr_696(8) or sumr_696(9));
E(326)<=not ( sumr_697(0) or sumr_697(1) or sumr_697(2) or sumr_697(3) or sumr_697(4) or sumr_697(5) or sumr_697(6) or sumr_697(7) or sumr_697(8) or sumr_697(9));
E(325)<=not ( sumr_698(0) or sumr_698(1) or sumr_698(2) or sumr_698(3) or sumr_698(4) or sumr_698(5) or sumr_698(6) or sumr_698(7) or sumr_698(8) or sumr_698(9));
E(324)<=not ( sumr_699(0) or sumr_699(1) or sumr_699(2) or sumr_699(3) or sumr_699(4) or sumr_699(5) or sumr_699(6) or sumr_699(7) or sumr_699(8) or sumr_699(9));
E(323)<=not ( sumr_700(0) or sumr_700(1) or sumr_700(2) or sumr_700(3) or sumr_700(4) or sumr_700(5) or sumr_700(6) or sumr_700(7) or sumr_700(8) or sumr_700(9));
E(322)<=not ( sumr_701(0) or sumr_701(1) or sumr_701(2) or sumr_701(3) or sumr_701(4) or sumr_701(5) or sumr_701(6) or sumr_701(7) or sumr_701(8) or sumr_701(9));
E(321)<=not ( sumr_702(0) or sumr_702(1) or sumr_702(2) or sumr_702(3) or sumr_702(4) or sumr_702(5) or sumr_702(6) or sumr_702(7) or sumr_702(8) or sumr_702(9));
E(320)<=not ( sumr_703(0) or sumr_703(1) or sumr_703(2) or sumr_703(3) or sumr_703(4) or sumr_703(5) or sumr_703(6) or sumr_703(7) or sumr_703(8) or sumr_703(9));
E(319)<=not ( sumr_704(0) or sumr_704(1) or sumr_704(2) or sumr_704(3) or sumr_704(4) or sumr_704(5) or sumr_704(6) or sumr_704(7) or sumr_704(8) or sumr_704(9));
E(318)<=not ( sumr_705(0) or sumr_705(1) or sumr_705(2) or sumr_705(3) or sumr_705(4) or sumr_705(5) or sumr_705(6) or sumr_705(7) or sumr_705(8) or sumr_705(9));
E(317)<=not ( sumr_706(0) or sumr_706(1) or sumr_706(2) or sumr_706(3) or sumr_706(4) or sumr_706(5) or sumr_706(6) or sumr_706(7) or sumr_706(8) or sumr_706(9));
E(316)<=not ( sumr_707(0) or sumr_707(1) or sumr_707(2) or sumr_707(3) or sumr_707(4) or sumr_707(5) or sumr_707(6) or sumr_707(7) or sumr_707(8) or sumr_707(9));
E(315)<=not ( sumr_708(0) or sumr_708(1) or sumr_708(2) or sumr_708(3) or sumr_708(4) or sumr_708(5) or sumr_708(6) or sumr_708(7) or sumr_708(8) or sumr_708(9));
E(314)<=not ( sumr_709(0) or sumr_709(1) or sumr_709(2) or sumr_709(3) or sumr_709(4) or sumr_709(5) or sumr_709(6) or sumr_709(7) or sumr_709(8) or sumr_709(9));
E(313)<=not ( sumr_710(0) or sumr_710(1) or sumr_710(2) or sumr_710(3) or sumr_710(4) or sumr_710(5) or sumr_710(6) or sumr_710(7) or sumr_710(8) or sumr_710(9));
E(312)<=not ( sumr_711(0) or sumr_711(1) or sumr_711(2) or sumr_711(3) or sumr_711(4) or sumr_711(5) or sumr_711(6) or sumr_711(7) or sumr_711(8) or sumr_711(9));
E(311)<=not ( sumr_712(0) or sumr_712(1) or sumr_712(2) or sumr_712(3) or sumr_712(4) or sumr_712(5) or sumr_712(6) or sumr_712(7) or sumr_712(8) or sumr_712(9));
E(310)<=not ( sumr_713(0) or sumr_713(1) or sumr_713(2) or sumr_713(3) or sumr_713(4) or sumr_713(5) or sumr_713(6) or sumr_713(7) or sumr_713(8) or sumr_713(9));
E(309)<=not ( sumr_714(0) or sumr_714(1) or sumr_714(2) or sumr_714(3) or sumr_714(4) or sumr_714(5) or sumr_714(6) or sumr_714(7) or sumr_714(8) or sumr_714(9));
E(308)<=not ( sumr_715(0) or sumr_715(1) or sumr_715(2) or sumr_715(3) or sumr_715(4) or sumr_715(5) or sumr_715(6) or sumr_715(7) or sumr_715(8) or sumr_715(9));
E(307)<=not ( sumr_716(0) or sumr_716(1) or sumr_716(2) or sumr_716(3) or sumr_716(4) or sumr_716(5) or sumr_716(6) or sumr_716(7) or sumr_716(8) or sumr_716(9));
E(306)<=not ( sumr_717(0) or sumr_717(1) or sumr_717(2) or sumr_717(3) or sumr_717(4) or sumr_717(5) or sumr_717(6) or sumr_717(7) or sumr_717(8) or sumr_717(9));
E(305)<=not ( sumr_718(0) or sumr_718(1) or sumr_718(2) or sumr_718(3) or sumr_718(4) or sumr_718(5) or sumr_718(6) or sumr_718(7) or sumr_718(8) or sumr_718(9));
E(304)<=not ( sumr_719(0) or sumr_719(1) or sumr_719(2) or sumr_719(3) or sumr_719(4) or sumr_719(5) or sumr_719(6) or sumr_719(7) or sumr_719(8) or sumr_719(9));
E(303)<=not ( sumr_720(0) or sumr_720(1) or sumr_720(2) or sumr_720(3) or sumr_720(4) or sumr_720(5) or sumr_720(6) or sumr_720(7) or sumr_720(8) or sumr_720(9));
E(302)<=not ( sumr_721(0) or sumr_721(1) or sumr_721(2) or sumr_721(3) or sumr_721(4) or sumr_721(5) or sumr_721(6) or sumr_721(7) or sumr_721(8) or sumr_721(9));
E(301)<=not ( sumr_722(0) or sumr_722(1) or sumr_722(2) or sumr_722(3) or sumr_722(4) or sumr_722(5) or sumr_722(6) or sumr_722(7) or sumr_722(8) or sumr_722(9));
E(300)<=not ( sumr_723(0) or sumr_723(1) or sumr_723(2) or sumr_723(3) or sumr_723(4) or sumr_723(5) or sumr_723(6) or sumr_723(7) or sumr_723(8) or sumr_723(9));
E(299)<=not ( sumr_724(0) or sumr_724(1) or sumr_724(2) or sumr_724(3) or sumr_724(4) or sumr_724(5) or sumr_724(6) or sumr_724(7) or sumr_724(8) or sumr_724(9));
E(298)<=not ( sumr_725(0) or sumr_725(1) or sumr_725(2) or sumr_725(3) or sumr_725(4) or sumr_725(5) or sumr_725(6) or sumr_725(7) or sumr_725(8) or sumr_725(9));
E(297)<=not ( sumr_726(0) or sumr_726(1) or sumr_726(2) or sumr_726(3) or sumr_726(4) or sumr_726(5) or sumr_726(6) or sumr_726(7) or sumr_726(8) or sumr_726(9));
E(296)<=not ( sumr_727(0) or sumr_727(1) or sumr_727(2) or sumr_727(3) or sumr_727(4) or sumr_727(5) or sumr_727(6) or sumr_727(7) or sumr_727(8) or sumr_727(9));
E(295)<=not ( sumr_728(0) or sumr_728(1) or sumr_728(2) or sumr_728(3) or sumr_728(4) or sumr_728(5) or sumr_728(6) or sumr_728(7) or sumr_728(8) or sumr_728(9));
E(294)<=not ( sumr_729(0) or sumr_729(1) or sumr_729(2) or sumr_729(3) or sumr_729(4) or sumr_729(5) or sumr_729(6) or sumr_729(7) or sumr_729(8) or sumr_729(9));
E(293)<=not ( sumr_730(0) or sumr_730(1) or sumr_730(2) or sumr_730(3) or sumr_730(4) or sumr_730(5) or sumr_730(6) or sumr_730(7) or sumr_730(8) or sumr_730(9));
E(292)<=not ( sumr_731(0) or sumr_731(1) or sumr_731(2) or sumr_731(3) or sumr_731(4) or sumr_731(5) or sumr_731(6) or sumr_731(7) or sumr_731(8) or sumr_731(9));
E(291)<=not ( sumr_732(0) or sumr_732(1) or sumr_732(2) or sumr_732(3) or sumr_732(4) or sumr_732(5) or sumr_732(6) or sumr_732(7) or sumr_732(8) or sumr_732(9));
E(290)<=not ( sumr_733(0) or sumr_733(1) or sumr_733(2) or sumr_733(3) or sumr_733(4) or sumr_733(5) or sumr_733(6) or sumr_733(7) or sumr_733(8) or sumr_733(9));
E(289)<=not ( sumr_734(0) or sumr_734(1) or sumr_734(2) or sumr_734(3) or sumr_734(4) or sumr_734(5) or sumr_734(6) or sumr_734(7) or sumr_734(8) or sumr_734(9));
E(288)<=not ( sumr_735(0) or sumr_735(1) or sumr_735(2) or sumr_735(3) or sumr_735(4) or sumr_735(5) or sumr_735(6) or sumr_735(7) or sumr_735(8) or sumr_735(9));
E(287)<=not ( sumr_736(0) or sumr_736(1) or sumr_736(2) or sumr_736(3) or sumr_736(4) or sumr_736(5) or sumr_736(6) or sumr_736(7) or sumr_736(8) or sumr_736(9));
E(286)<=not ( sumr_737(0) or sumr_737(1) or sumr_737(2) or sumr_737(3) or sumr_737(4) or sumr_737(5) or sumr_737(6) or sumr_737(7) or sumr_737(8) or sumr_737(9));
E(285)<=not ( sumr_738(0) or sumr_738(1) or sumr_738(2) or sumr_738(3) or sumr_738(4) or sumr_738(5) or sumr_738(6) or sumr_738(7) or sumr_738(8) or sumr_738(9));
E(284)<=not ( sumr_739(0) or sumr_739(1) or sumr_739(2) or sumr_739(3) or sumr_739(4) or sumr_739(5) or sumr_739(6) or sumr_739(7) or sumr_739(8) or sumr_739(9));
E(283)<=not ( sumr_740(0) or sumr_740(1) or sumr_740(2) or sumr_740(3) or sumr_740(4) or sumr_740(5) or sumr_740(6) or sumr_740(7) or sumr_740(8) or sumr_740(9));
E(282)<=not ( sumr_741(0) or sumr_741(1) or sumr_741(2) or sumr_741(3) or sumr_741(4) or sumr_741(5) or sumr_741(6) or sumr_741(7) or sumr_741(8) or sumr_741(9));
E(281)<=not ( sumr_742(0) or sumr_742(1) or sumr_742(2) or sumr_742(3) or sumr_742(4) or sumr_742(5) or sumr_742(6) or sumr_742(7) or sumr_742(8) or sumr_742(9));
E(280)<=not ( sumr_743(0) or sumr_743(1) or sumr_743(2) or sumr_743(3) or sumr_743(4) or sumr_743(5) or sumr_743(6) or sumr_743(7) or sumr_743(8) or sumr_743(9));
E(279)<=not ( sumr_744(0) or sumr_744(1) or sumr_744(2) or sumr_744(3) or sumr_744(4) or sumr_744(5) or sumr_744(6) or sumr_744(7) or sumr_744(8) or sumr_744(9));
E(278)<=not ( sumr_745(0) or sumr_745(1) or sumr_745(2) or sumr_745(3) or sumr_745(4) or sumr_745(5) or sumr_745(6) or sumr_745(7) or sumr_745(8) or sumr_745(9));
E(277)<=not ( sumr_746(0) or sumr_746(1) or sumr_746(2) or sumr_746(3) or sumr_746(4) or sumr_746(5) or sumr_746(6) or sumr_746(7) or sumr_746(8) or sumr_746(9));
E(276)<=not ( sumr_747(0) or sumr_747(1) or sumr_747(2) or sumr_747(3) or sumr_747(4) or sumr_747(5) or sumr_747(6) or sumr_747(7) or sumr_747(8) or sumr_747(9));
E(275)<=not ( sumr_748(0) or sumr_748(1) or sumr_748(2) or sumr_748(3) or sumr_748(4) or sumr_748(5) or sumr_748(6) or sumr_748(7) or sumr_748(8) or sumr_748(9));
E(274)<=not ( sumr_749(0) or sumr_749(1) or sumr_749(2) or sumr_749(3) or sumr_749(4) or sumr_749(5) or sumr_749(6) or sumr_749(7) or sumr_749(8) or sumr_749(9));
E(273)<=not ( sumr_750(0) or sumr_750(1) or sumr_750(2) or sumr_750(3) or sumr_750(4) or sumr_750(5) or sumr_750(6) or sumr_750(7) or sumr_750(8) or sumr_750(9));
E(272)<=not ( sumr_751(0) or sumr_751(1) or sumr_751(2) or sumr_751(3) or sumr_751(4) or sumr_751(5) or sumr_751(6) or sumr_751(7) or sumr_751(8) or sumr_751(9));
E(271)<=not ( sumr_752(0) or sumr_752(1) or sumr_752(2) or sumr_752(3) or sumr_752(4) or sumr_752(5) or sumr_752(6) or sumr_752(7) or sumr_752(8) or sumr_752(9));
E(270)<=not ( sumr_753(0) or sumr_753(1) or sumr_753(2) or sumr_753(3) or sumr_753(4) or sumr_753(5) or sumr_753(6) or sumr_753(7) or sumr_753(8) or sumr_753(9));
E(269)<=not ( sumr_754(0) or sumr_754(1) or sumr_754(2) or sumr_754(3) or sumr_754(4) or sumr_754(5) or sumr_754(6) or sumr_754(7) or sumr_754(8) or sumr_754(9));
E(268)<=not ( sumr_755(0) or sumr_755(1) or sumr_755(2) or sumr_755(3) or sumr_755(4) or sumr_755(5) or sumr_755(6) or sumr_755(7) or sumr_755(8) or sumr_755(9));
E(267)<=not ( sumr_756(0) or sumr_756(1) or sumr_756(2) or sumr_756(3) or sumr_756(4) or sumr_756(5) or sumr_756(6) or sumr_756(7) or sumr_756(8) or sumr_756(9));
E(266)<=not ( sumr_757(0) or sumr_757(1) or sumr_757(2) or sumr_757(3) or sumr_757(4) or sumr_757(5) or sumr_757(6) or sumr_757(7) or sumr_757(8) or sumr_757(9));
E(265)<=not ( sumr_758(0) or sumr_758(1) or sumr_758(2) or sumr_758(3) or sumr_758(4) or sumr_758(5) or sumr_758(6) or sumr_758(7) or sumr_758(8) or sumr_758(9));
E(264)<=not ( sumr_759(0) or sumr_759(1) or sumr_759(2) or sumr_759(3) or sumr_759(4) or sumr_759(5) or sumr_759(6) or sumr_759(7) or sumr_759(8) or sumr_759(9));
E(263)<=not ( sumr_760(0) or sumr_760(1) or sumr_760(2) or sumr_760(3) or sumr_760(4) or sumr_760(5) or sumr_760(6) or sumr_760(7) or sumr_760(8) or sumr_760(9));
E(262)<=not ( sumr_761(0) or sumr_761(1) or sumr_761(2) or sumr_761(3) or sumr_761(4) or sumr_761(5) or sumr_761(6) or sumr_761(7) or sumr_761(8) or sumr_761(9));
E(261)<=not ( sumr_762(0) or sumr_762(1) or sumr_762(2) or sumr_762(3) or sumr_762(4) or sumr_762(5) or sumr_762(6) or sumr_762(7) or sumr_762(8) or sumr_762(9));
E(260)<=not ( sumr_763(0) or sumr_763(1) or sumr_763(2) or sumr_763(3) or sumr_763(4) or sumr_763(5) or sumr_763(6) or sumr_763(7) or sumr_763(8) or sumr_763(9));
E(259)<=not ( sumr_764(0) or sumr_764(1) or sumr_764(2) or sumr_764(3) or sumr_764(4) or sumr_764(5) or sumr_764(6) or sumr_764(7) or sumr_764(8) or sumr_764(9));
E(258)<=not ( sumr_765(0) or sumr_765(1) or sumr_765(2) or sumr_765(3) or sumr_765(4) or sumr_765(5) or sumr_765(6) or sumr_765(7) or sumr_765(8) or sumr_765(9));
E(257)<=not ( sumr_766(0) or sumr_766(1) or sumr_766(2) or sumr_766(3) or sumr_766(4) or sumr_766(5) or sumr_766(6) or sumr_766(7) or sumr_766(8) or sumr_766(9));
E(256)<=not ( sumr_767(0) or sumr_767(1) or sumr_767(2) or sumr_767(3) or sumr_767(4) or sumr_767(5) or sumr_767(6) or sumr_767(7) or sumr_767(8) or sumr_767(9));
E(255)<=not ( sumr_768(0) or sumr_768(1) or sumr_768(2) or sumr_768(3) or sumr_768(4) or sumr_768(5) or sumr_768(6) or sumr_768(7) or sumr_768(8) or sumr_768(9));
E(254)<=not ( sumr_769(0) or sumr_769(1) or sumr_769(2) or sumr_769(3) or sumr_769(4) or sumr_769(5) or sumr_769(6) or sumr_769(7) or sumr_769(8) or sumr_769(9));
E(253)<=not ( sumr_770(0) or sumr_770(1) or sumr_770(2) or sumr_770(3) or sumr_770(4) or sumr_770(5) or sumr_770(6) or sumr_770(7) or sumr_770(8) or sumr_770(9));
E(252)<=not ( sumr_771(0) or sumr_771(1) or sumr_771(2) or sumr_771(3) or sumr_771(4) or sumr_771(5) or sumr_771(6) or sumr_771(7) or sumr_771(8) or sumr_771(9));
E(251)<=not ( sumr_772(0) or sumr_772(1) or sumr_772(2) or sumr_772(3) or sumr_772(4) or sumr_772(5) or sumr_772(6) or sumr_772(7) or sumr_772(8) or sumr_772(9));
E(250)<=not ( sumr_773(0) or sumr_773(1) or sumr_773(2) or sumr_773(3) or sumr_773(4) or sumr_773(5) or sumr_773(6) or sumr_773(7) or sumr_773(8) or sumr_773(9));
E(249)<=not ( sumr_774(0) or sumr_774(1) or sumr_774(2) or sumr_774(3) or sumr_774(4) or sumr_774(5) or sumr_774(6) or sumr_774(7) or sumr_774(8) or sumr_774(9));
E(248)<=not ( sumr_775(0) or sumr_775(1) or sumr_775(2) or sumr_775(3) or sumr_775(4) or sumr_775(5) or sumr_775(6) or sumr_775(7) or sumr_775(8) or sumr_775(9));
E(247)<=not ( sumr_776(0) or sumr_776(1) or sumr_776(2) or sumr_776(3) or sumr_776(4) or sumr_776(5) or sumr_776(6) or sumr_776(7) or sumr_776(8) or sumr_776(9));
E(246)<=not ( sumr_777(0) or sumr_777(1) or sumr_777(2) or sumr_777(3) or sumr_777(4) or sumr_777(5) or sumr_777(6) or sumr_777(7) or sumr_777(8) or sumr_777(9));
E(245)<=not ( sumr_778(0) or sumr_778(1) or sumr_778(2) or sumr_778(3) or sumr_778(4) or sumr_778(5) or sumr_778(6) or sumr_778(7) or sumr_778(8) or sumr_778(9));
E(244)<=not ( sumr_779(0) or sumr_779(1) or sumr_779(2) or sumr_779(3) or sumr_779(4) or sumr_779(5) or sumr_779(6) or sumr_779(7) or sumr_779(8) or sumr_779(9));
E(243)<=not ( sumr_780(0) or sumr_780(1) or sumr_780(2) or sumr_780(3) or sumr_780(4) or sumr_780(5) or sumr_780(6) or sumr_780(7) or sumr_780(8) or sumr_780(9));
E(242)<=not ( sumr_781(0) or sumr_781(1) or sumr_781(2) or sumr_781(3) or sumr_781(4) or sumr_781(5) or sumr_781(6) or sumr_781(7) or sumr_781(8) or sumr_781(9));
E(241)<=not ( sumr_782(0) or sumr_782(1) or sumr_782(2) or sumr_782(3) or sumr_782(4) or sumr_782(5) or sumr_782(6) or sumr_782(7) or sumr_782(8) or sumr_782(9));
E(240)<=not ( sumr_783(0) or sumr_783(1) or sumr_783(2) or sumr_783(3) or sumr_783(4) or sumr_783(5) or sumr_783(6) or sumr_783(7) or sumr_783(8) or sumr_783(9));
E(239)<=not ( sumr_784(0) or sumr_784(1) or sumr_784(2) or sumr_784(3) or sumr_784(4) or sumr_784(5) or sumr_784(6) or sumr_784(7) or sumr_784(8) or sumr_784(9));
E(238)<=not ( sumr_785(0) or sumr_785(1) or sumr_785(2) or sumr_785(3) or sumr_785(4) or sumr_785(5) or sumr_785(6) or sumr_785(7) or sumr_785(8) or sumr_785(9));
E(237)<=not ( sumr_786(0) or sumr_786(1) or sumr_786(2) or sumr_786(3) or sumr_786(4) or sumr_786(5) or sumr_786(6) or sumr_786(7) or sumr_786(8) or sumr_786(9));
E(236)<=not ( sumr_787(0) or sumr_787(1) or sumr_787(2) or sumr_787(3) or sumr_787(4) or sumr_787(5) or sumr_787(6) or sumr_787(7) or sumr_787(8) or sumr_787(9));
E(235)<=not ( sumr_788(0) or sumr_788(1) or sumr_788(2) or sumr_788(3) or sumr_788(4) or sumr_788(5) or sumr_788(6) or sumr_788(7) or sumr_788(8) or sumr_788(9));
E(234)<=not ( sumr_789(0) or sumr_789(1) or sumr_789(2) or sumr_789(3) or sumr_789(4) or sumr_789(5) or sumr_789(6) or sumr_789(7) or sumr_789(8) or sumr_789(9));
E(233)<=not ( sumr_790(0) or sumr_790(1) or sumr_790(2) or sumr_790(3) or sumr_790(4) or sumr_790(5) or sumr_790(6) or sumr_790(7) or sumr_790(8) or sumr_790(9));
E(232)<=not ( sumr_791(0) or sumr_791(1) or sumr_791(2) or sumr_791(3) or sumr_791(4) or sumr_791(5) or sumr_791(6) or sumr_791(7) or sumr_791(8) or sumr_791(9));
E(231)<=not ( sumr_792(0) or sumr_792(1) or sumr_792(2) or sumr_792(3) or sumr_792(4) or sumr_792(5) or sumr_792(6) or sumr_792(7) or sumr_792(8) or sumr_792(9));
E(230)<=not ( sumr_793(0) or sumr_793(1) or sumr_793(2) or sumr_793(3) or sumr_793(4) or sumr_793(5) or sumr_793(6) or sumr_793(7) or sumr_793(8) or sumr_793(9));
E(229)<=not ( sumr_794(0) or sumr_794(1) or sumr_794(2) or sumr_794(3) or sumr_794(4) or sumr_794(5) or sumr_794(6) or sumr_794(7) or sumr_794(8) or sumr_794(9));
E(228)<=not ( sumr_795(0) or sumr_795(1) or sumr_795(2) or sumr_795(3) or sumr_795(4) or sumr_795(5) or sumr_795(6) or sumr_795(7) or sumr_795(8) or sumr_795(9));
E(227)<=not ( sumr_796(0) or sumr_796(1) or sumr_796(2) or sumr_796(3) or sumr_796(4) or sumr_796(5) or sumr_796(6) or sumr_796(7) or sumr_796(8) or sumr_796(9));
E(226)<=not ( sumr_797(0) or sumr_797(1) or sumr_797(2) or sumr_797(3) or sumr_797(4) or sumr_797(5) or sumr_797(6) or sumr_797(7) or sumr_797(8) or sumr_797(9));
E(225)<=not ( sumr_798(0) or sumr_798(1) or sumr_798(2) or sumr_798(3) or sumr_798(4) or sumr_798(5) or sumr_798(6) or sumr_798(7) or sumr_798(8) or sumr_798(9));
E(224)<=not ( sumr_799(0) or sumr_799(1) or sumr_799(2) or sumr_799(3) or sumr_799(4) or sumr_799(5) or sumr_799(6) or sumr_799(7) or sumr_799(8) or sumr_799(9));
E(223)<=not ( sumr_800(0) or sumr_800(1) or sumr_800(2) or sumr_800(3) or sumr_800(4) or sumr_800(5) or sumr_800(6) or sumr_800(7) or sumr_800(8) or sumr_800(9));
E(222)<=not ( sumr_801(0) or sumr_801(1) or sumr_801(2) or sumr_801(3) or sumr_801(4) or sumr_801(5) or sumr_801(6) or sumr_801(7) or sumr_801(8) or sumr_801(9));
E(221)<=not ( sumr_802(0) or sumr_802(1) or sumr_802(2) or sumr_802(3) or sumr_802(4) or sumr_802(5) or sumr_802(6) or sumr_802(7) or sumr_802(8) or sumr_802(9));
E(220)<=not ( sumr_803(0) or sumr_803(1) or sumr_803(2) or sumr_803(3) or sumr_803(4) or sumr_803(5) or sumr_803(6) or sumr_803(7) or sumr_803(8) or sumr_803(9));
E(219)<=not ( sumr_804(0) or sumr_804(1) or sumr_804(2) or sumr_804(3) or sumr_804(4) or sumr_804(5) or sumr_804(6) or sumr_804(7) or sumr_804(8) or sumr_804(9));
E(218)<=not ( sumr_805(0) or sumr_805(1) or sumr_805(2) or sumr_805(3) or sumr_805(4) or sumr_805(5) or sumr_805(6) or sumr_805(7) or sumr_805(8) or sumr_805(9));
E(217)<=not ( sumr_806(0) or sumr_806(1) or sumr_806(2) or sumr_806(3) or sumr_806(4) or sumr_806(5) or sumr_806(6) or sumr_806(7) or sumr_806(8) or sumr_806(9));
E(216)<=not ( sumr_807(0) or sumr_807(1) or sumr_807(2) or sumr_807(3) or sumr_807(4) or sumr_807(5) or sumr_807(6) or sumr_807(7) or sumr_807(8) or sumr_807(9));
E(215)<=not ( sumr_808(0) or sumr_808(1) or sumr_808(2) or sumr_808(3) or sumr_808(4) or sumr_808(5) or sumr_808(6) or sumr_808(7) or sumr_808(8) or sumr_808(9));
E(214)<=not ( sumr_809(0) or sumr_809(1) or sumr_809(2) or sumr_809(3) or sumr_809(4) or sumr_809(5) or sumr_809(6) or sumr_809(7) or sumr_809(8) or sumr_809(9));
E(213)<=not ( sumr_810(0) or sumr_810(1) or sumr_810(2) or sumr_810(3) or sumr_810(4) or sumr_810(5) or sumr_810(6) or sumr_810(7) or sumr_810(8) or sumr_810(9));
E(212)<=not ( sumr_811(0) or sumr_811(1) or sumr_811(2) or sumr_811(3) or sumr_811(4) or sumr_811(5) or sumr_811(6) or sumr_811(7) or sumr_811(8) or sumr_811(9));
E(211)<=not ( sumr_812(0) or sumr_812(1) or sumr_812(2) or sumr_812(3) or sumr_812(4) or sumr_812(5) or sumr_812(6) or sumr_812(7) or sumr_812(8) or sumr_812(9));
E(210)<=not ( sumr_813(0) or sumr_813(1) or sumr_813(2) or sumr_813(3) or sumr_813(4) or sumr_813(5) or sumr_813(6) or sumr_813(7) or sumr_813(8) or sumr_813(9));
E(209)<=not ( sumr_814(0) or sumr_814(1) or sumr_814(2) or sumr_814(3) or sumr_814(4) or sumr_814(5) or sumr_814(6) or sumr_814(7) or sumr_814(8) or sumr_814(9));
E(208)<=not ( sumr_815(0) or sumr_815(1) or sumr_815(2) or sumr_815(3) or sumr_815(4) or sumr_815(5) or sumr_815(6) or sumr_815(7) or sumr_815(8) or sumr_815(9));
E(207)<=not ( sumr_816(0) or sumr_816(1) or sumr_816(2) or sumr_816(3) or sumr_816(4) or sumr_816(5) or sumr_816(6) or sumr_816(7) or sumr_816(8) or sumr_816(9));
E(206)<=not ( sumr_817(0) or sumr_817(1) or sumr_817(2) or sumr_817(3) or sumr_817(4) or sumr_817(5) or sumr_817(6) or sumr_817(7) or sumr_817(8) or sumr_817(9));
E(205)<=not ( sumr_818(0) or sumr_818(1) or sumr_818(2) or sumr_818(3) or sumr_818(4) or sumr_818(5) or sumr_818(6) or sumr_818(7) or sumr_818(8) or sumr_818(9));
E(204)<=not ( sumr_819(0) or sumr_819(1) or sumr_819(2) or sumr_819(3) or sumr_819(4) or sumr_819(5) or sumr_819(6) or sumr_819(7) or sumr_819(8) or sumr_819(9));
E(203)<=not ( sumr_820(0) or sumr_820(1) or sumr_820(2) or sumr_820(3) or sumr_820(4) or sumr_820(5) or sumr_820(6) or sumr_820(7) or sumr_820(8) or sumr_820(9));
E(202)<=not ( sumr_821(0) or sumr_821(1) or sumr_821(2) or sumr_821(3) or sumr_821(4) or sumr_821(5) or sumr_821(6) or sumr_821(7) or sumr_821(8) or sumr_821(9));
E(201)<=not ( sumr_822(0) or sumr_822(1) or sumr_822(2) or sumr_822(3) or sumr_822(4) or sumr_822(5) or sumr_822(6) or sumr_822(7) or sumr_822(8) or sumr_822(9));
E(200)<=not ( sumr_823(0) or sumr_823(1) or sumr_823(2) or sumr_823(3) or sumr_823(4) or sumr_823(5) or sumr_823(6) or sumr_823(7) or sumr_823(8) or sumr_823(9));
E(199)<=not ( sumr_824(0) or sumr_824(1) or sumr_824(2) or sumr_824(3) or sumr_824(4) or sumr_824(5) or sumr_824(6) or sumr_824(7) or sumr_824(8) or sumr_824(9));
E(198)<=not ( sumr_825(0) or sumr_825(1) or sumr_825(2) or sumr_825(3) or sumr_825(4) or sumr_825(5) or sumr_825(6) or sumr_825(7) or sumr_825(8) or sumr_825(9));
E(197)<=not ( sumr_826(0) or sumr_826(1) or sumr_826(2) or sumr_826(3) or sumr_826(4) or sumr_826(5) or sumr_826(6) or sumr_826(7) or sumr_826(8) or sumr_826(9));
E(196)<=not ( sumr_827(0) or sumr_827(1) or sumr_827(2) or sumr_827(3) or sumr_827(4) or sumr_827(5) or sumr_827(6) or sumr_827(7) or sumr_827(8) or sumr_827(9));
E(195)<=not ( sumr_828(0) or sumr_828(1) or sumr_828(2) or sumr_828(3) or sumr_828(4) or sumr_828(5) or sumr_828(6) or sumr_828(7) or sumr_828(8) or sumr_828(9));
E(194)<=not ( sumr_829(0) or sumr_829(1) or sumr_829(2) or sumr_829(3) or sumr_829(4) or sumr_829(5) or sumr_829(6) or sumr_829(7) or sumr_829(8) or sumr_829(9));
E(193)<=not ( sumr_830(0) or sumr_830(1) or sumr_830(2) or sumr_830(3) or sumr_830(4) or sumr_830(5) or sumr_830(6) or sumr_830(7) or sumr_830(8) or sumr_830(9));
E(192)<=not ( sumr_831(0) or sumr_831(1) or sumr_831(2) or sumr_831(3) or sumr_831(4) or sumr_831(5) or sumr_831(6) or sumr_831(7) or sumr_831(8) or sumr_831(9));
E(191)<=not ( sumr_832(0) or sumr_832(1) or sumr_832(2) or sumr_832(3) or sumr_832(4) or sumr_832(5) or sumr_832(6) or sumr_832(7) or sumr_832(8) or sumr_832(9));
E(190)<=not ( sumr_833(0) or sumr_833(1) or sumr_833(2) or sumr_833(3) or sumr_833(4) or sumr_833(5) or sumr_833(6) or sumr_833(7) or sumr_833(8) or sumr_833(9));
E(189)<=not ( sumr_834(0) or sumr_834(1) or sumr_834(2) or sumr_834(3) or sumr_834(4) or sumr_834(5) or sumr_834(6) or sumr_834(7) or sumr_834(8) or sumr_834(9));
E(188)<=not ( sumr_835(0) or sumr_835(1) or sumr_835(2) or sumr_835(3) or sumr_835(4) or sumr_835(5) or sumr_835(6) or sumr_835(7) or sumr_835(8) or sumr_835(9));
E(187)<=not ( sumr_836(0) or sumr_836(1) or sumr_836(2) or sumr_836(3) or sumr_836(4) or sumr_836(5) or sumr_836(6) or sumr_836(7) or sumr_836(8) or sumr_836(9));
E(186)<=not ( sumr_837(0) or sumr_837(1) or sumr_837(2) or sumr_837(3) or sumr_837(4) or sumr_837(5) or sumr_837(6) or sumr_837(7) or sumr_837(8) or sumr_837(9));
E(185)<=not ( sumr_838(0) or sumr_838(1) or sumr_838(2) or sumr_838(3) or sumr_838(4) or sumr_838(5) or sumr_838(6) or sumr_838(7) or sumr_838(8) or sumr_838(9));
E(184)<=not ( sumr_839(0) or sumr_839(1) or sumr_839(2) or sumr_839(3) or sumr_839(4) or sumr_839(5) or sumr_839(6) or sumr_839(7) or sumr_839(8) or sumr_839(9));
E(183)<=not ( sumr_840(0) or sumr_840(1) or sumr_840(2) or sumr_840(3) or sumr_840(4) or sumr_840(5) or sumr_840(6) or sumr_840(7) or sumr_840(8) or sumr_840(9));
E(182)<=not ( sumr_841(0) or sumr_841(1) or sumr_841(2) or sumr_841(3) or sumr_841(4) or sumr_841(5) or sumr_841(6) or sumr_841(7) or sumr_841(8) or sumr_841(9));
E(181)<=not ( sumr_842(0) or sumr_842(1) or sumr_842(2) or sumr_842(3) or sumr_842(4) or sumr_842(5) or sumr_842(6) or sumr_842(7) or sumr_842(8) or sumr_842(9));
E(180)<=not ( sumr_843(0) or sumr_843(1) or sumr_843(2) or sumr_843(3) or sumr_843(4) or sumr_843(5) or sumr_843(6) or sumr_843(7) or sumr_843(8) or sumr_843(9));
E(179)<=not ( sumr_844(0) or sumr_844(1) or sumr_844(2) or sumr_844(3) or sumr_844(4) or sumr_844(5) or sumr_844(6) or sumr_844(7) or sumr_844(8) or sumr_844(9));
E(178)<=not ( sumr_845(0) or sumr_845(1) or sumr_845(2) or sumr_845(3) or sumr_845(4) or sumr_845(5) or sumr_845(6) or sumr_845(7) or sumr_845(8) or sumr_845(9));
E(177)<=not ( sumr_846(0) or sumr_846(1) or sumr_846(2) or sumr_846(3) or sumr_846(4) or sumr_846(5) or sumr_846(6) or sumr_846(7) or sumr_846(8) or sumr_846(9));
E(176)<=not ( sumr_847(0) or sumr_847(1) or sumr_847(2) or sumr_847(3) or sumr_847(4) or sumr_847(5) or sumr_847(6) or sumr_847(7) or sumr_847(8) or sumr_847(9));
E(175)<=not ( sumr_848(0) or sumr_848(1) or sumr_848(2) or sumr_848(3) or sumr_848(4) or sumr_848(5) or sumr_848(6) or sumr_848(7) or sumr_848(8) or sumr_848(9));
E(174)<=not ( sumr_849(0) or sumr_849(1) or sumr_849(2) or sumr_849(3) or sumr_849(4) or sumr_849(5) or sumr_849(6) or sumr_849(7) or sumr_849(8) or sumr_849(9));
E(173)<=not ( sumr_850(0) or sumr_850(1) or sumr_850(2) or sumr_850(3) or sumr_850(4) or sumr_850(5) or sumr_850(6) or sumr_850(7) or sumr_850(8) or sumr_850(9));
E(172)<=not ( sumr_851(0) or sumr_851(1) or sumr_851(2) or sumr_851(3) or sumr_851(4) or sumr_851(5) or sumr_851(6) or sumr_851(7) or sumr_851(8) or sumr_851(9));
E(171)<=not ( sumr_852(0) or sumr_852(1) or sumr_852(2) or sumr_852(3) or sumr_852(4) or sumr_852(5) or sumr_852(6) or sumr_852(7) or sumr_852(8) or sumr_852(9));
E(170)<=not ( sumr_853(0) or sumr_853(1) or sumr_853(2) or sumr_853(3) or sumr_853(4) or sumr_853(5) or sumr_853(6) or sumr_853(7) or sumr_853(8) or sumr_853(9));
E(169)<=not ( sumr_854(0) or sumr_854(1) or sumr_854(2) or sumr_854(3) or sumr_854(4) or sumr_854(5) or sumr_854(6) or sumr_854(7) or sumr_854(8) or sumr_854(9));
E(168)<=not ( sumr_855(0) or sumr_855(1) or sumr_855(2) or sumr_855(3) or sumr_855(4) or sumr_855(5) or sumr_855(6) or sumr_855(7) or sumr_855(8) or sumr_855(9));
E(167)<=not ( sumr_856(0) or sumr_856(1) or sumr_856(2) or sumr_856(3) or sumr_856(4) or sumr_856(5) or sumr_856(6) or sumr_856(7) or sumr_856(8) or sumr_856(9));
E(166)<=not ( sumr_857(0) or sumr_857(1) or sumr_857(2) or sumr_857(3) or sumr_857(4) or sumr_857(5) or sumr_857(6) or sumr_857(7) or sumr_857(8) or sumr_857(9));
E(165)<=not ( sumr_858(0) or sumr_858(1) or sumr_858(2) or sumr_858(3) or sumr_858(4) or sumr_858(5) or sumr_858(6) or sumr_858(7) or sumr_858(8) or sumr_858(9));
E(164)<=not ( sumr_859(0) or sumr_859(1) or sumr_859(2) or sumr_859(3) or sumr_859(4) or sumr_859(5) or sumr_859(6) or sumr_859(7) or sumr_859(8) or sumr_859(9));
E(163)<=not ( sumr_860(0) or sumr_860(1) or sumr_860(2) or sumr_860(3) or sumr_860(4) or sumr_860(5) or sumr_860(6) or sumr_860(7) or sumr_860(8) or sumr_860(9));
E(162)<=not ( sumr_861(0) or sumr_861(1) or sumr_861(2) or sumr_861(3) or sumr_861(4) or sumr_861(5) or sumr_861(6) or sumr_861(7) or sumr_861(8) or sumr_861(9));
E(161)<=not ( sumr_862(0) or sumr_862(1) or sumr_862(2) or sumr_862(3) or sumr_862(4) or sumr_862(5) or sumr_862(6) or sumr_862(7) or sumr_862(8) or sumr_862(9));
E(160)<=not ( sumr_863(0) or sumr_863(1) or sumr_863(2) or sumr_863(3) or sumr_863(4) or sumr_863(5) or sumr_863(6) or sumr_863(7) or sumr_863(8) or sumr_863(9));
E(159)<=not ( sumr_864(0) or sumr_864(1) or sumr_864(2) or sumr_864(3) or sumr_864(4) or sumr_864(5) or sumr_864(6) or sumr_864(7) or sumr_864(8) or sumr_864(9));
E(158)<=not ( sumr_865(0) or sumr_865(1) or sumr_865(2) or sumr_865(3) or sumr_865(4) or sumr_865(5) or sumr_865(6) or sumr_865(7) or sumr_865(8) or sumr_865(9));
E(157)<=not ( sumr_866(0) or sumr_866(1) or sumr_866(2) or sumr_866(3) or sumr_866(4) or sumr_866(5) or sumr_866(6) or sumr_866(7) or sumr_866(8) or sumr_866(9));
E(156)<=not ( sumr_867(0) or sumr_867(1) or sumr_867(2) or sumr_867(3) or sumr_867(4) or sumr_867(5) or sumr_867(6) or sumr_867(7) or sumr_867(8) or sumr_867(9));
E(155)<=not ( sumr_868(0) or sumr_868(1) or sumr_868(2) or sumr_868(3) or sumr_868(4) or sumr_868(5) or sumr_868(6) or sumr_868(7) or sumr_868(8) or sumr_868(9));
E(154)<=not ( sumr_869(0) or sumr_869(1) or sumr_869(2) or sumr_869(3) or sumr_869(4) or sumr_869(5) or sumr_869(6) or sumr_869(7) or sumr_869(8) or sumr_869(9));
E(153)<=not ( sumr_870(0) or sumr_870(1) or sumr_870(2) or sumr_870(3) or sumr_870(4) or sumr_870(5) or sumr_870(6) or sumr_870(7) or sumr_870(8) or sumr_870(9));
E(152)<=not ( sumr_871(0) or sumr_871(1) or sumr_871(2) or sumr_871(3) or sumr_871(4) or sumr_871(5) or sumr_871(6) or sumr_871(7) or sumr_871(8) or sumr_871(9));
E(151)<=not ( sumr_872(0) or sumr_872(1) or sumr_872(2) or sumr_872(3) or sumr_872(4) or sumr_872(5) or sumr_872(6) or sumr_872(7) or sumr_872(8) or sumr_872(9));
E(150)<=not ( sumr_873(0) or sumr_873(1) or sumr_873(2) or sumr_873(3) or sumr_873(4) or sumr_873(5) or sumr_873(6) or sumr_873(7) or sumr_873(8) or sumr_873(9));
E(149)<=not ( sumr_874(0) or sumr_874(1) or sumr_874(2) or sumr_874(3) or sumr_874(4) or sumr_874(5) or sumr_874(6) or sumr_874(7) or sumr_874(8) or sumr_874(9));
E(148)<=not ( sumr_875(0) or sumr_875(1) or sumr_875(2) or sumr_875(3) or sumr_875(4) or sumr_875(5) or sumr_875(6) or sumr_875(7) or sumr_875(8) or sumr_875(9));
E(147)<=not ( sumr_876(0) or sumr_876(1) or sumr_876(2) or sumr_876(3) or sumr_876(4) or sumr_876(5) or sumr_876(6) or sumr_876(7) or sumr_876(8) or sumr_876(9));
E(146)<=not ( sumr_877(0) or sumr_877(1) or sumr_877(2) or sumr_877(3) or sumr_877(4) or sumr_877(5) or sumr_877(6) or sumr_877(7) or sumr_877(8) or sumr_877(9));
E(145)<=not ( sumr_878(0) or sumr_878(1) or sumr_878(2) or sumr_878(3) or sumr_878(4) or sumr_878(5) or sumr_878(6) or sumr_878(7) or sumr_878(8) or sumr_878(9));
E(144)<=not ( sumr_879(0) or sumr_879(1) or sumr_879(2) or sumr_879(3) or sumr_879(4) or sumr_879(5) or sumr_879(6) or sumr_879(7) or sumr_879(8) or sumr_879(9));
E(143)<=not ( sumr_880(0) or sumr_880(1) or sumr_880(2) or sumr_880(3) or sumr_880(4) or sumr_880(5) or sumr_880(6) or sumr_880(7) or sumr_880(8) or sumr_880(9));
E(142)<=not ( sumr_881(0) or sumr_881(1) or sumr_881(2) or sumr_881(3) or sumr_881(4) or sumr_881(5) or sumr_881(6) or sumr_881(7) or sumr_881(8) or sumr_881(9));
E(141)<=not ( sumr_882(0) or sumr_882(1) or sumr_882(2) or sumr_882(3) or sumr_882(4) or sumr_882(5) or sumr_882(6) or sumr_882(7) or sumr_882(8) or sumr_882(9));
E(140)<=not ( sumr_883(0) or sumr_883(1) or sumr_883(2) or sumr_883(3) or sumr_883(4) or sumr_883(5) or sumr_883(6) or sumr_883(7) or sumr_883(8) or sumr_883(9));
E(139)<=not ( sumr_884(0) or sumr_884(1) or sumr_884(2) or sumr_884(3) or sumr_884(4) or sumr_884(5) or sumr_884(6) or sumr_884(7) or sumr_884(8) or sumr_884(9));
E(138)<=not ( sumr_885(0) or sumr_885(1) or sumr_885(2) or sumr_885(3) or sumr_885(4) or sumr_885(5) or sumr_885(6) or sumr_885(7) or sumr_885(8) or sumr_885(9));
E(137)<=not ( sumr_886(0) or sumr_886(1) or sumr_886(2) or sumr_886(3) or sumr_886(4) or sumr_886(5) or sumr_886(6) or sumr_886(7) or sumr_886(8) or sumr_886(9));
E(136)<=not ( sumr_887(0) or sumr_887(1) or sumr_887(2) or sumr_887(3) or sumr_887(4) or sumr_887(5) or sumr_887(6) or sumr_887(7) or sumr_887(8) or sumr_887(9));
E(135)<=not ( sumr_888(0) or sumr_888(1) or sumr_888(2) or sumr_888(3) or sumr_888(4) or sumr_888(5) or sumr_888(6) or sumr_888(7) or sumr_888(8) or sumr_888(9));
E(134)<=not ( sumr_889(0) or sumr_889(1) or sumr_889(2) or sumr_889(3) or sumr_889(4) or sumr_889(5) or sumr_889(6) or sumr_889(7) or sumr_889(8) or sumr_889(9));
E(133)<=not ( sumr_890(0) or sumr_890(1) or sumr_890(2) or sumr_890(3) or sumr_890(4) or sumr_890(5) or sumr_890(6) or sumr_890(7) or sumr_890(8) or sumr_890(9));
E(132)<=not ( sumr_891(0) or sumr_891(1) or sumr_891(2) or sumr_891(3) or sumr_891(4) or sumr_891(5) or sumr_891(6) or sumr_891(7) or sumr_891(8) or sumr_891(9));
E(131)<=not ( sumr_892(0) or sumr_892(1) or sumr_892(2) or sumr_892(3) or sumr_892(4) or sumr_892(5) or sumr_892(6) or sumr_892(7) or sumr_892(8) or sumr_892(9));
E(130)<=not ( sumr_893(0) or sumr_893(1) or sumr_893(2) or sumr_893(3) or sumr_893(4) or sumr_893(5) or sumr_893(6) or sumr_893(7) or sumr_893(8) or sumr_893(9));
E(129)<=not ( sumr_894(0) or sumr_894(1) or sumr_894(2) or sumr_894(3) or sumr_894(4) or sumr_894(5) or sumr_894(6) or sumr_894(7) or sumr_894(8) or sumr_894(9));
E(128)<=not ( sumr_895(0) or sumr_895(1) or sumr_895(2) or sumr_895(3) or sumr_895(4) or sumr_895(5) or sumr_895(6) or sumr_895(7) or sumr_895(8) or sumr_895(9));
E(127)<=not ( sumr_896(0) or sumr_896(1) or sumr_896(2) or sumr_896(3) or sumr_896(4) or sumr_896(5) or sumr_896(6) or sumr_896(7) or sumr_896(8) or sumr_896(9));
E(126)<=not ( sumr_897(0) or sumr_897(1) or sumr_897(2) or sumr_897(3) or sumr_897(4) or sumr_897(5) or sumr_897(6) or sumr_897(7) or sumr_897(8) or sumr_897(9));
E(125)<=not ( sumr_898(0) or sumr_898(1) or sumr_898(2) or sumr_898(3) or sumr_898(4) or sumr_898(5) or sumr_898(6) or sumr_898(7) or sumr_898(8) or sumr_898(9));
E(124)<=not ( sumr_899(0) or sumr_899(1) or sumr_899(2) or sumr_899(3) or sumr_899(4) or sumr_899(5) or sumr_899(6) or sumr_899(7) or sumr_899(8) or sumr_899(9));
E(123)<=not ( sumr_900(0) or sumr_900(1) or sumr_900(2) or sumr_900(3) or sumr_900(4) or sumr_900(5) or sumr_900(6) or sumr_900(7) or sumr_900(8) or sumr_900(9));
E(122)<=not ( sumr_901(0) or sumr_901(1) or sumr_901(2) or sumr_901(3) or sumr_901(4) or sumr_901(5) or sumr_901(6) or sumr_901(7) or sumr_901(8) or sumr_901(9));
E(121)<=not ( sumr_902(0) or sumr_902(1) or sumr_902(2) or sumr_902(3) or sumr_902(4) or sumr_902(5) or sumr_902(6) or sumr_902(7) or sumr_902(8) or sumr_902(9));
E(120)<=not ( sumr_903(0) or sumr_903(1) or sumr_903(2) or sumr_903(3) or sumr_903(4) or sumr_903(5) or sumr_903(6) or sumr_903(7) or sumr_903(8) or sumr_903(9));
E(119)<=not ( sumr_904(0) or sumr_904(1) or sumr_904(2) or sumr_904(3) or sumr_904(4) or sumr_904(5) or sumr_904(6) or sumr_904(7) or sumr_904(8) or sumr_904(9));
E(118)<=not ( sumr_905(0) or sumr_905(1) or sumr_905(2) or sumr_905(3) or sumr_905(4) or sumr_905(5) or sumr_905(6) or sumr_905(7) or sumr_905(8) or sumr_905(9));
E(117)<=not ( sumr_906(0) or sumr_906(1) or sumr_906(2) or sumr_906(3) or sumr_906(4) or sumr_906(5) or sumr_906(6) or sumr_906(7) or sumr_906(8) or sumr_906(9));
E(116)<=not ( sumr_907(0) or sumr_907(1) or sumr_907(2) or sumr_907(3) or sumr_907(4) or sumr_907(5) or sumr_907(6) or sumr_907(7) or sumr_907(8) or sumr_907(9));
E(115)<=not ( sumr_908(0) or sumr_908(1) or sumr_908(2) or sumr_908(3) or sumr_908(4) or sumr_908(5) or sumr_908(6) or sumr_908(7) or sumr_908(8) or sumr_908(9));
E(114)<=not ( sumr_909(0) or sumr_909(1) or sumr_909(2) or sumr_909(3) or sumr_909(4) or sumr_909(5) or sumr_909(6) or sumr_909(7) or sumr_909(8) or sumr_909(9));
E(113)<=not ( sumr_910(0) or sumr_910(1) or sumr_910(2) or sumr_910(3) or sumr_910(4) or sumr_910(5) or sumr_910(6) or sumr_910(7) or sumr_910(8) or sumr_910(9));
E(112)<=not ( sumr_911(0) or sumr_911(1) or sumr_911(2) or sumr_911(3) or sumr_911(4) or sumr_911(5) or sumr_911(6) or sumr_911(7) or sumr_911(8) or sumr_911(9));
E(111)<=not ( sumr_912(0) or sumr_912(1) or sumr_912(2) or sumr_912(3) or sumr_912(4) or sumr_912(5) or sumr_912(6) or sumr_912(7) or sumr_912(8) or sumr_912(9));
E(110)<=not ( sumr_913(0) or sumr_913(1) or sumr_913(2) or sumr_913(3) or sumr_913(4) or sumr_913(5) or sumr_913(6) or sumr_913(7) or sumr_913(8) or sumr_913(9));
E(109)<=not ( sumr_914(0) or sumr_914(1) or sumr_914(2) or sumr_914(3) or sumr_914(4) or sumr_914(5) or sumr_914(6) or sumr_914(7) or sumr_914(8) or sumr_914(9));
E(108)<=not ( sumr_915(0) or sumr_915(1) or sumr_915(2) or sumr_915(3) or sumr_915(4) or sumr_915(5) or sumr_915(6) or sumr_915(7) or sumr_915(8) or sumr_915(9));
E(107)<=not ( sumr_916(0) or sumr_916(1) or sumr_916(2) or sumr_916(3) or sumr_916(4) or sumr_916(5) or sumr_916(6) or sumr_916(7) or sumr_916(8) or sumr_916(9));
E(106)<=not ( sumr_917(0) or sumr_917(1) or sumr_917(2) or sumr_917(3) or sumr_917(4) or sumr_917(5) or sumr_917(6) or sumr_917(7) or sumr_917(8) or sumr_917(9));
E(105)<=not ( sumr_918(0) or sumr_918(1) or sumr_918(2) or sumr_918(3) or sumr_918(4) or sumr_918(5) or sumr_918(6) or sumr_918(7) or sumr_918(8) or sumr_918(9));
E(104)<=not ( sumr_919(0) or sumr_919(1) or sumr_919(2) or sumr_919(3) or sumr_919(4) or sumr_919(5) or sumr_919(6) or sumr_919(7) or sumr_919(8) or sumr_919(9));
E(103)<=not ( sumr_920(0) or sumr_920(1) or sumr_920(2) or sumr_920(3) or sumr_920(4) or sumr_920(5) or sumr_920(6) or sumr_920(7) or sumr_920(8) or sumr_920(9));
E(102)<=not ( sumr_921(0) or sumr_921(1) or sumr_921(2) or sumr_921(3) or sumr_921(4) or sumr_921(5) or sumr_921(6) or sumr_921(7) or sumr_921(8) or sumr_921(9));
E(101)<=not ( sumr_922(0) or sumr_922(1) or sumr_922(2) or sumr_922(3) or sumr_922(4) or sumr_922(5) or sumr_922(6) or sumr_922(7) or sumr_922(8) or sumr_922(9));
E(100)<=not ( sumr_923(0) or sumr_923(1) or sumr_923(2) or sumr_923(3) or sumr_923(4) or sumr_923(5) or sumr_923(6) or sumr_923(7) or sumr_923(8) or sumr_923(9));
E(99)<=not ( sumr_924(0) or sumr_924(1) or sumr_924(2) or sumr_924(3) or sumr_924(4) or sumr_924(5) or sumr_924(6) or sumr_924(7) or sumr_924(8) or sumr_924(9));
E(98)<=not ( sumr_925(0) or sumr_925(1) or sumr_925(2) or sumr_925(3) or sumr_925(4) or sumr_925(5) or sumr_925(6) or sumr_925(7) or sumr_925(8) or sumr_925(9));
E(97)<=not ( sumr_926(0) or sumr_926(1) or sumr_926(2) or sumr_926(3) or sumr_926(4) or sumr_926(5) or sumr_926(6) or sumr_926(7) or sumr_926(8) or sumr_926(9));
E(96)<=not ( sumr_927(0) or sumr_927(1) or sumr_927(2) or sumr_927(3) or sumr_927(4) or sumr_927(5) or sumr_927(6) or sumr_927(7) or sumr_927(8) or sumr_927(9));
E(95)<=not ( sumr_928(0) or sumr_928(1) or sumr_928(2) or sumr_928(3) or sumr_928(4) or sumr_928(5) or sumr_928(6) or sumr_928(7) or sumr_928(8) or sumr_928(9));
E(94)<=not ( sumr_929(0) or sumr_929(1) or sumr_929(2) or sumr_929(3) or sumr_929(4) or sumr_929(5) or sumr_929(6) or sumr_929(7) or sumr_929(8) or sumr_929(9));
E(93)<=not ( sumr_930(0) or sumr_930(1) or sumr_930(2) or sumr_930(3) or sumr_930(4) or sumr_930(5) or sumr_930(6) or sumr_930(7) or sumr_930(8) or sumr_930(9));
E(92)<=not ( sumr_931(0) or sumr_931(1) or sumr_931(2) or sumr_931(3) or sumr_931(4) or sumr_931(5) or sumr_931(6) or sumr_931(7) or sumr_931(8) or sumr_931(9));
E(91)<=not ( sumr_932(0) or sumr_932(1) or sumr_932(2) or sumr_932(3) or sumr_932(4) or sumr_932(5) or sumr_932(6) or sumr_932(7) or sumr_932(8) or sumr_932(9));
E(90)<=not ( sumr_933(0) or sumr_933(1) or sumr_933(2) or sumr_933(3) or sumr_933(4) or sumr_933(5) or sumr_933(6) or sumr_933(7) or sumr_933(8) or sumr_933(9));
E(89)<=not ( sumr_934(0) or sumr_934(1) or sumr_934(2) or sumr_934(3) or sumr_934(4) or sumr_934(5) or sumr_934(6) or sumr_934(7) or sumr_934(8) or sumr_934(9));
E(88)<=not ( sumr_935(0) or sumr_935(1) or sumr_935(2) or sumr_935(3) or sumr_935(4) or sumr_935(5) or sumr_935(6) or sumr_935(7) or sumr_935(8) or sumr_935(9));
E(87)<=not ( sumr_936(0) or sumr_936(1) or sumr_936(2) or sumr_936(3) or sumr_936(4) or sumr_936(5) or sumr_936(6) or sumr_936(7) or sumr_936(8) or sumr_936(9));
E(86)<=not ( sumr_937(0) or sumr_937(1) or sumr_937(2) or sumr_937(3) or sumr_937(4) or sumr_937(5) or sumr_937(6) or sumr_937(7) or sumr_937(8) or sumr_937(9));
E(85)<=not ( sumr_938(0) or sumr_938(1) or sumr_938(2) or sumr_938(3) or sumr_938(4) or sumr_938(5) or sumr_938(6) or sumr_938(7) or sumr_938(8) or sumr_938(9));
E(84)<=not ( sumr_939(0) or sumr_939(1) or sumr_939(2) or sumr_939(3) or sumr_939(4) or sumr_939(5) or sumr_939(6) or sumr_939(7) or sumr_939(8) or sumr_939(9));
E(83)<=not ( sumr_940(0) or sumr_940(1) or sumr_940(2) or sumr_940(3) or sumr_940(4) or sumr_940(5) or sumr_940(6) or sumr_940(7) or sumr_940(8) or sumr_940(9));
E(82)<=not ( sumr_941(0) or sumr_941(1) or sumr_941(2) or sumr_941(3) or sumr_941(4) or sumr_941(5) or sumr_941(6) or sumr_941(7) or sumr_941(8) or sumr_941(9));
E(81)<=not ( sumr_942(0) or sumr_942(1) or sumr_942(2) or sumr_942(3) or sumr_942(4) or sumr_942(5) or sumr_942(6) or sumr_942(7) or sumr_942(8) or sumr_942(9));
E(80)<=not ( sumr_943(0) or sumr_943(1) or sumr_943(2) or sumr_943(3) or sumr_943(4) or sumr_943(5) or sumr_943(6) or sumr_943(7) or sumr_943(8) or sumr_943(9));
E(79)<=not ( sumr_944(0) or sumr_944(1) or sumr_944(2) or sumr_944(3) or sumr_944(4) or sumr_944(5) or sumr_944(6) or sumr_944(7) or sumr_944(8) or sumr_944(9));
E(78)<=not ( sumr_945(0) or sumr_945(1) or sumr_945(2) or sumr_945(3) or sumr_945(4) or sumr_945(5) or sumr_945(6) or sumr_945(7) or sumr_945(8) or sumr_945(9));
E(77)<=not ( sumr_946(0) or sumr_946(1) or sumr_946(2) or sumr_946(3) or sumr_946(4) or sumr_946(5) or sumr_946(6) or sumr_946(7) or sumr_946(8) or sumr_946(9));
E(76)<=not ( sumr_947(0) or sumr_947(1) or sumr_947(2) or sumr_947(3) or sumr_947(4) or sumr_947(5) or sumr_947(6) or sumr_947(7) or sumr_947(8) or sumr_947(9));
E(75)<=not ( sumr_948(0) or sumr_948(1) or sumr_948(2) or sumr_948(3) or sumr_948(4) or sumr_948(5) or sumr_948(6) or sumr_948(7) or sumr_948(8) or sumr_948(9));
E(74)<=not ( sumr_949(0) or sumr_949(1) or sumr_949(2) or sumr_949(3) or sumr_949(4) or sumr_949(5) or sumr_949(6) or sumr_949(7) or sumr_949(8) or sumr_949(9));
E(73)<=not ( sumr_950(0) or sumr_950(1) or sumr_950(2) or sumr_950(3) or sumr_950(4) or sumr_950(5) or sumr_950(6) or sumr_950(7) or sumr_950(8) or sumr_950(9));
E(72)<=not ( sumr_951(0) or sumr_951(1) or sumr_951(2) or sumr_951(3) or sumr_951(4) or sumr_951(5) or sumr_951(6) or sumr_951(7) or sumr_951(8) or sumr_951(9));
E(71)<=not ( sumr_952(0) or sumr_952(1) or sumr_952(2) or sumr_952(3) or sumr_952(4) or sumr_952(5) or sumr_952(6) or sumr_952(7) or sumr_952(8) or sumr_952(9));
E(70)<=not ( sumr_953(0) or sumr_953(1) or sumr_953(2) or sumr_953(3) or sumr_953(4) or sumr_953(5) or sumr_953(6) or sumr_953(7) or sumr_953(8) or sumr_953(9));
E(69)<=not ( sumr_954(0) or sumr_954(1) or sumr_954(2) or sumr_954(3) or sumr_954(4) or sumr_954(5) or sumr_954(6) or sumr_954(7) or sumr_954(8) or sumr_954(9));
E(68)<=not ( sumr_955(0) or sumr_955(1) or sumr_955(2) or sumr_955(3) or sumr_955(4) or sumr_955(5) or sumr_955(6) or sumr_955(7) or sumr_955(8) or sumr_955(9));
E(67)<=not ( sumr_956(0) or sumr_956(1) or sumr_956(2) or sumr_956(3) or sumr_956(4) or sumr_956(5) or sumr_956(6) or sumr_956(7) or sumr_956(8) or sumr_956(9));
E(66)<=not ( sumr_957(0) or sumr_957(1) or sumr_957(2) or sumr_957(3) or sumr_957(4) or sumr_957(5) or sumr_957(6) or sumr_957(7) or sumr_957(8) or sumr_957(9));
E(65)<=not ( sumr_958(0) or sumr_958(1) or sumr_958(2) or sumr_958(3) or sumr_958(4) or sumr_958(5) or sumr_958(6) or sumr_958(7) or sumr_958(8) or sumr_958(9));
E(64)<=not ( sumr_959(0) or sumr_959(1) or sumr_959(2) or sumr_959(3) or sumr_959(4) or sumr_959(5) or sumr_959(6) or sumr_959(7) or sumr_959(8) or sumr_959(9));
E(63)<=not ( sumr_960(0) or sumr_960(1) or sumr_960(2) or sumr_960(3) or sumr_960(4) or sumr_960(5) or sumr_960(6) or sumr_960(7) or sumr_960(8) or sumr_960(9));
E(62)<=not ( sumr_961(0) or sumr_961(1) or sumr_961(2) or sumr_961(3) or sumr_961(4) or sumr_961(5) or sumr_961(6) or sumr_961(7) or sumr_961(8) or sumr_961(9));
E(61)<=not ( sumr_962(0) or sumr_962(1) or sumr_962(2) or sumr_962(3) or sumr_962(4) or sumr_962(5) or sumr_962(6) or sumr_962(7) or sumr_962(8) or sumr_962(9));
E(60)<=not ( sumr_963(0) or sumr_963(1) or sumr_963(2) or sumr_963(3) or sumr_963(4) or sumr_963(5) or sumr_963(6) or sumr_963(7) or sumr_963(8) or sumr_963(9));
E(59)<=not ( sumr_964(0) or sumr_964(1) or sumr_964(2) or sumr_964(3) or sumr_964(4) or sumr_964(5) or sumr_964(6) or sumr_964(7) or sumr_964(8) or sumr_964(9));
E(58)<=not ( sumr_965(0) or sumr_965(1) or sumr_965(2) or sumr_965(3) or sumr_965(4) or sumr_965(5) or sumr_965(6) or sumr_965(7) or sumr_965(8) or sumr_965(9));
E(57)<=not ( sumr_966(0) or sumr_966(1) or sumr_966(2) or sumr_966(3) or sumr_966(4) or sumr_966(5) or sumr_966(6) or sumr_966(7) or sumr_966(8) or sumr_966(9));
E(56)<=not ( sumr_967(0) or sumr_967(1) or sumr_967(2) or sumr_967(3) or sumr_967(4) or sumr_967(5) or sumr_967(6) or sumr_967(7) or sumr_967(8) or sumr_967(9));
E(55)<=not ( sumr_968(0) or sumr_968(1) or sumr_968(2) or sumr_968(3) or sumr_968(4) or sumr_968(5) or sumr_968(6) or sumr_968(7) or sumr_968(8) or sumr_968(9));
E(54)<=not ( sumr_969(0) or sumr_969(1) or sumr_969(2) or sumr_969(3) or sumr_969(4) or sumr_969(5) or sumr_969(6) or sumr_969(7) or sumr_969(8) or sumr_969(9));
E(53)<=not ( sumr_970(0) or sumr_970(1) or sumr_970(2) or sumr_970(3) or sumr_970(4) or sumr_970(5) or sumr_970(6) or sumr_970(7) or sumr_970(8) or sumr_970(9));
E(52)<=not ( sumr_971(0) or sumr_971(1) or sumr_971(2) or sumr_971(3) or sumr_971(4) or sumr_971(5) or sumr_971(6) or sumr_971(7) or sumr_971(8) or sumr_971(9));
E(51)<=not ( sumr_972(0) or sumr_972(1) or sumr_972(2) or sumr_972(3) or sumr_972(4) or sumr_972(5) or sumr_972(6) or sumr_972(7) or sumr_972(8) or sumr_972(9));
E(50)<=not ( sumr_973(0) or sumr_973(1) or sumr_973(2) or sumr_973(3) or sumr_973(4) or sumr_973(5) or sumr_973(6) or sumr_973(7) or sumr_973(8) or sumr_973(9));
E(49)<=not ( sumr_974(0) or sumr_974(1) or sumr_974(2) or sumr_974(3) or sumr_974(4) or sumr_974(5) or sumr_974(6) or sumr_974(7) or sumr_974(8) or sumr_974(9));
E(48)<=not ( sumr_975(0) or sumr_975(1) or sumr_975(2) or sumr_975(3) or sumr_975(4) or sumr_975(5) or sumr_975(6) or sumr_975(7) or sumr_975(8) or sumr_975(9));
E(47)<=not ( sumr_976(0) or sumr_976(1) or sumr_976(2) or sumr_976(3) or sumr_976(4) or sumr_976(5) or sumr_976(6) or sumr_976(7) or sumr_976(8) or sumr_976(9));
E(46)<=not ( sumr_977(0) or sumr_977(1) or sumr_977(2) or sumr_977(3) or sumr_977(4) or sumr_977(5) or sumr_977(6) or sumr_977(7) or sumr_977(8) or sumr_977(9));
E(45)<=not ( sumr_978(0) or sumr_978(1) or sumr_978(2) or sumr_978(3) or sumr_978(4) or sumr_978(5) or sumr_978(6) or sumr_978(7) or sumr_978(8) or sumr_978(9));
E(44)<=not ( sumr_979(0) or sumr_979(1) or sumr_979(2) or sumr_979(3) or sumr_979(4) or sumr_979(5) or sumr_979(6) or sumr_979(7) or sumr_979(8) or sumr_979(9));
E(43)<=not ( sumr_980(0) or sumr_980(1) or sumr_980(2) or sumr_980(3) or sumr_980(4) or sumr_980(5) or sumr_980(6) or sumr_980(7) or sumr_980(8) or sumr_980(9));
E(42)<=not ( sumr_981(0) or sumr_981(1) or sumr_981(2) or sumr_981(3) or sumr_981(4) or sumr_981(5) or sumr_981(6) or sumr_981(7) or sumr_981(8) or sumr_981(9));
E(41)<=not ( sumr_982(0) or sumr_982(1) or sumr_982(2) or sumr_982(3) or sumr_982(4) or sumr_982(5) or sumr_982(6) or sumr_982(7) or sumr_982(8) or sumr_982(9));
E(40)<=not ( sumr_983(0) or sumr_983(1) or sumr_983(2) or sumr_983(3) or sumr_983(4) or sumr_983(5) or sumr_983(6) or sumr_983(7) or sumr_983(8) or sumr_983(9));
E(39)<=not ( sumr_984(0) or sumr_984(1) or sumr_984(2) or sumr_984(3) or sumr_984(4) or sumr_984(5) or sumr_984(6) or sumr_984(7) or sumr_984(8) or sumr_984(9));
E(38)<=not ( sumr_985(0) or sumr_985(1) or sumr_985(2) or sumr_985(3) or sumr_985(4) or sumr_985(5) or sumr_985(6) or sumr_985(7) or sumr_985(8) or sumr_985(9));
E(37)<=not ( sumr_986(0) or sumr_986(1) or sumr_986(2) or sumr_986(3) or sumr_986(4) or sumr_986(5) or sumr_986(6) or sumr_986(7) or sumr_986(8) or sumr_986(9));
E(36)<=not ( sumr_987(0) or sumr_987(1) or sumr_987(2) or sumr_987(3) or sumr_987(4) or sumr_987(5) or sumr_987(6) or sumr_987(7) or sumr_987(8) or sumr_987(9));
E(35)<=not ( sumr_988(0) or sumr_988(1) or sumr_988(2) or sumr_988(3) or sumr_988(4) or sumr_988(5) or sumr_988(6) or sumr_988(7) or sumr_988(8) or sumr_988(9));
E(34)<=not ( sumr_989(0) or sumr_989(1) or sumr_989(2) or sumr_989(3) or sumr_989(4) or sumr_989(5) or sumr_989(6) or sumr_989(7) or sumr_989(8) or sumr_989(9));
E(33)<=not ( sumr_990(0) or sumr_990(1) or sumr_990(2) or sumr_990(3) or sumr_990(4) or sumr_990(5) or sumr_990(6) or sumr_990(7) or sumr_990(8) or sumr_990(9));
E(32)<=not ( sumr_991(0) or sumr_991(1) or sumr_991(2) or sumr_991(3) or sumr_991(4) or sumr_991(5) or sumr_991(6) or sumr_991(7) or sumr_991(8) or sumr_991(9));
E(31)<=not ( sumr_992(0) or sumr_992(1) or sumr_992(2) or sumr_992(3) or sumr_992(4) or sumr_992(5) or sumr_992(6) or sumr_992(7) or sumr_992(8) or sumr_992(9));
E(30)<=not ( sumr_993(0) or sumr_993(1) or sumr_993(2) or sumr_993(3) or sumr_993(4) or sumr_993(5) or sumr_993(6) or sumr_993(7) or sumr_993(8) or sumr_993(9));
E(29)<=not ( sumr_994(0) or sumr_994(1) or sumr_994(2) or sumr_994(3) or sumr_994(4) or sumr_994(5) or sumr_994(6) or sumr_994(7) or sumr_994(8) or sumr_994(9));
E(28)<=not ( sumr_995(0) or sumr_995(1) or sumr_995(2) or sumr_995(3) or sumr_995(4) or sumr_995(5) or sumr_995(6) or sumr_995(7) or sumr_995(8) or sumr_995(9));
E(27)<=not ( sumr_996(0) or sumr_996(1) or sumr_996(2) or sumr_996(3) or sumr_996(4) or sumr_996(5) or sumr_996(6) or sumr_996(7) or sumr_996(8) or sumr_996(9));
E(26)<=not ( sumr_997(0) or sumr_997(1) or sumr_997(2) or sumr_997(3) or sumr_997(4) or sumr_997(5) or sumr_997(6) or sumr_997(7) or sumr_997(8) or sumr_997(9));
E(25)<=not ( sumr_998(0) or sumr_998(1) or sumr_998(2) or sumr_998(3) or sumr_998(4) or sumr_998(5) or sumr_998(6) or sumr_998(7) or sumr_998(8) or sumr_998(9));
E(24)<=not ( sumr_999(0) or sumr_999(1) or sumr_999(2) or sumr_999(3) or sumr_999(4) or sumr_999(5) or sumr_999(6) or sumr_999(7) or sumr_999(8) or sumr_999(9));
E(23)<=not ( sumr_1000(0) or sumr_1000(1) or sumr_1000(2) or sumr_1000(3) or sumr_1000(4) or sumr_1000(5) or sumr_1000(6) or sumr_1000(7) or sumr_1000(8) or sumr_1000(9));
E(22)<=not ( sumr_1001(0) or sumr_1001(1) or sumr_1001(2) or sumr_1001(3) or sumr_1001(4) or sumr_1001(5) or sumr_1001(6) or sumr_1001(7) or sumr_1001(8) or sumr_1001(9));
E(21)<=not ( sumr_1002(0) or sumr_1002(1) or sumr_1002(2) or sumr_1002(3) or sumr_1002(4) or sumr_1002(5) or sumr_1002(6) or sumr_1002(7) or sumr_1002(8) or sumr_1002(9));
E(20)<=not ( sumr_1003(0) or sumr_1003(1) or sumr_1003(2) or sumr_1003(3) or sumr_1003(4) or sumr_1003(5) or sumr_1003(6) or sumr_1003(7) or sumr_1003(8) or sumr_1003(9));
E(19)<=not ( sumr_1004(0) or sumr_1004(1) or sumr_1004(2) or sumr_1004(3) or sumr_1004(4) or sumr_1004(5) or sumr_1004(6) or sumr_1004(7) or sumr_1004(8) or sumr_1004(9));
E(18)<=not ( sumr_1005(0) or sumr_1005(1) or sumr_1005(2) or sumr_1005(3) or sumr_1005(4) or sumr_1005(5) or sumr_1005(6) or sumr_1005(7) or sumr_1005(8) or sumr_1005(9));
E(17)<=not ( sumr_1006(0) or sumr_1006(1) or sumr_1006(2) or sumr_1006(3) or sumr_1006(4) or sumr_1006(5) or sumr_1006(6) or sumr_1006(7) or sumr_1006(8) or sumr_1006(9));
E(16)<=not ( sumr_1007(0) or sumr_1007(1) or sumr_1007(2) or sumr_1007(3) or sumr_1007(4) or sumr_1007(5) or sumr_1007(6) or sumr_1007(7) or sumr_1007(8) or sumr_1007(9));
E(15)<=not ( sumr_1008(0) or sumr_1008(1) or sumr_1008(2) or sumr_1008(3) or sumr_1008(4) or sumr_1008(5) or sumr_1008(6) or sumr_1008(7) or sumr_1008(8) or sumr_1008(9));
E(14)<=not ( sumr_1009(0) or sumr_1009(1) or sumr_1009(2) or sumr_1009(3) or sumr_1009(4) or sumr_1009(5) or sumr_1009(6) or sumr_1009(7) or sumr_1009(8) or sumr_1009(9));
E(13)<=not ( sumr_1010(0) or sumr_1010(1) or sumr_1010(2) or sumr_1010(3) or sumr_1010(4) or sumr_1010(5) or sumr_1010(6) or sumr_1010(7) or sumr_1010(8) or sumr_1010(9));
E(12)<=not ( sumr_1011(0) or sumr_1011(1) or sumr_1011(2) or sumr_1011(3) or sumr_1011(4) or sumr_1011(5) or sumr_1011(6) or sumr_1011(7) or sumr_1011(8) or sumr_1011(9));
E(11)<=not ( sumr_1012(0) or sumr_1012(1) or sumr_1012(2) or sumr_1012(3) or sumr_1012(4) or sumr_1012(5) or sumr_1012(6) or sumr_1012(7) or sumr_1012(8) or sumr_1012(9));
E(10)<=not ( sumr_1013(0) or sumr_1013(1) or sumr_1013(2) or sumr_1013(3) or sumr_1013(4) or sumr_1013(5) or sumr_1013(6) or sumr_1013(7) or sumr_1013(8) or sumr_1013(9));
E(9)<=not ( sumr_1014(0) or sumr_1014(1) or sumr_1014(2) or sumr_1014(3) or sumr_1014(4) or sumr_1014(5) or sumr_1014(6) or sumr_1014(7) or sumr_1014(8) or sumr_1014(9));
E(8)<=not ( sumr_1015(0) or sumr_1015(1) or sumr_1015(2) or sumr_1015(3) or sumr_1015(4) or sumr_1015(5) or sumr_1015(6) or sumr_1015(7) or sumr_1015(8) or sumr_1015(9));
E(7)<=not ( sumr_1016(0) or sumr_1016(1) or sumr_1016(2) or sumr_1016(3) or sumr_1016(4) or sumr_1016(5) or sumr_1016(6) or sumr_1016(7) or sumr_1016(8) or sumr_1016(9));
E(6)<=not ( sumr_1017(0) or sumr_1017(1) or sumr_1017(2) or sumr_1017(3) or sumr_1017(4) or sumr_1017(5) or sumr_1017(6) or sumr_1017(7) or sumr_1017(8) or sumr_1017(9));
E(5)<=not ( sumr_1018(0) or sumr_1018(1) or sumr_1018(2) or sumr_1018(3) or sumr_1018(4) or sumr_1018(5) or sumr_1018(6) or sumr_1018(7) or sumr_1018(8) or sumr_1018(9));
E(4)<=not ( sumr_1019(0) or sumr_1019(1) or sumr_1019(2) or sumr_1019(3) or sumr_1019(4) or sumr_1019(5) or sumr_1019(6) or sumr_1019(7) or sumr_1019(8) or sumr_1019(9));
E(3)<=not ( sumr_1020(0) or sumr_1020(1) or sumr_1020(2) or sumr_1020(3) or sumr_1020(4) or sumr_1020(5) or sumr_1020(6) or sumr_1020(7) or sumr_1020(8) or sumr_1020(9));
E(2)<=not ( sumr_1021(0) or sumr_1021(1) or sumr_1021(2) or sumr_1021(3) or sumr_1021(4) or sumr_1021(5) or sumr_1021(6) or sumr_1021(7) or sumr_1021(8) or sumr_1021(9));
E(1)<=not ( sumr_1022(0) or sumr_1022(1) or sumr_1022(2) or sumr_1022(3) or sumr_1022(4) or sumr_1022(5) or sumr_1022(6) or sumr_1022(7) or sumr_1022(8) or sumr_1022(9));
E(0)<=not ( sumr_1023(0) or sumr_1023(1) or sumr_1023(2) or sumr_1023(3) or sumr_1023(4) or sumr_1023(5) or sumr_1023(6) or sumr_1023(7) or sumr_1023(8) or sumr_1023(9));
end arch;
