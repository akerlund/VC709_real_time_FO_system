library ieee;
use ieee.std_logic_1164.all;
entity synenc is
    port(
        in_data     :    in  std_logic_vector(1012 downto 0);
        out_data    :    out std_logic_vector(1022 downto 0)
);
end entity;

architecture arch of synenc is
begin
out_data(1012 downto 0) <= in_data;
out_data(1022)<= in_data(1012) xor in_data(1009) xor in_data(1006) xor in_data(1003) xor in_data(1002) xor in_data(1000) xor in_data(997) xor in_data(996) xor in_data(994) xor in_data(992) xor in_data(991) xor in_data(990) xor in_data(989) xor in_data(988) xor in_data(985) xor in_data(984) xor in_data(980) xor in_data(979) xor in_data(978) xor in_data(977) xor in_data(976) xor in_data(973) xor in_data(969) xor in_data(968) xor in_data(967) xor in_data(965) xor in_data(964) xor in_data(963) xor in_data(962) xor in_data(961) xor in_data(960) xor in_data(955) xor in_data(954) xor in_data(953) xor in_data(945) xor in_data(944) xor in_data(943) xor in_data(942) xor in_data(941) xor in_data(940) xor in_data(939) xor in_data(938) xor in_data(937) xor in_data(936) xor in_data(932) xor in_data(931) xor in_data(930) xor in_data(926) xor in_data(923) xor in_data(922) xor in_data(921) xor in_data(919) xor in_data(918) xor in_data(915) xor in_data(913) xor in_data(911) xor in_data(910) xor in_data(909) xor in_data(907) xor in_data(906) xor in_data(905) xor in_data(904) xor in_data(902) xor in_data(900) xor in_data(896) xor in_data(895) xor in_data(894) xor in_data(893) xor in_data(891) xor in_data(888) xor in_data(886) xor in_data(884) xor in_data(878) xor in_data(876) xor in_data(875) xor in_data(874) xor in_data(873) xor in_data(872) xor in_data(871) xor in_data(870) xor in_data(869) xor in_data(867) xor in_data(865) xor in_data(863) xor in_data(861) xor in_data(859) xor in_data(858) xor in_data(857) xor in_data(856) xor in_data(854) xor in_data(849) xor in_data(848) xor in_data(847) xor in_data(845) xor in_data(842) xor in_data(838) xor in_data(837) xor in_data(834) xor in_data(832) xor in_data(831) xor in_data(829) xor in_data(827) xor in_data(826) xor in_data(823) xor in_data(822) xor in_data(821) xor in_data(820) xor in_data(818) xor in_data(816) xor in_data(815) xor in_data(811) xor in_data(810) xor in_data(807) xor in_data(806) xor in_data(805) xor in_data(804) xor in_data(803) xor in_data(802) xor in_data(799) xor in_data(797) xor in_data(795) xor in_data(793) xor in_data(790) xor in_data(789) xor in_data(786) xor in_data(785) xor in_data(782) xor in_data(780) xor in_data(777) xor in_data(776) xor in_data(775) xor in_data(774) xor in_data(773) xor in_data(771) xor in_data(768) xor in_data(767) xor in_data(766) xor in_data(761) xor in_data(757) xor in_data(756) xor in_data(754) xor in_data(753) xor in_data(750) xor in_data(746) xor in_data(744) xor in_data(741) xor in_data(740) xor in_data(738) xor in_data(737) xor in_data(736) xor in_data(735) xor in_data(733) xor in_data(732) xor in_data(731) xor in_data(729) xor in_data(727) xor in_data(725) xor in_data(724) xor in_data(723) xor in_data(720) xor in_data(719) xor in_data(716) xor in_data(715) xor in_data(714) xor in_data(712) xor in_data(711) xor in_data(710) xor in_data(708) xor in_data(707) xor in_data(706) xor in_data(703) xor in_data(702) xor in_data(701) xor in_data(699) xor in_data(697) xor in_data(694) xor in_data(693) xor in_data(692) xor in_data(690) xor in_data(684) xor in_data(683) xor in_data(682) xor in_data(681) xor in_data(679) xor in_data(678) xor in_data(676) xor in_data(675) xor in_data(674) xor in_data(669) xor in_data(668) xor in_data(664) xor in_data(661) xor in_data(659) xor in_data(656) xor in_data(654) xor in_data(653) xor in_data(650) xor in_data(649) xor in_data(647) xor in_data(643) xor in_data(639) xor in_data(637) xor in_data(636) xor in_data(634) xor in_data(631) xor in_data(629) xor in_data(628) xor in_data(627) xor in_data(625) xor in_data(622) xor in_data(621) xor in_data(617) xor in_data(615) xor in_data(614) xor in_data(607) xor in_data(605) xor in_data(602) xor in_data(599) xor in_data(597) xor in_data(596) xor in_data(595) xor in_data(594) xor in_data(593) xor in_data(591) xor in_data(590) xor in_data(589) xor in_data(588) xor in_data(584) xor in_data(583) xor in_data(579) xor in_data(578) xor in_data(576) xor in_data(575) xor in_data(574) xor in_data(572) xor in_data(571) xor in_data(566) xor in_data(565) xor in_data(564) xor in_data(563) xor in_data(560) xor in_data(557) xor in_data(556) xor in_data(555) xor in_data(552) xor in_data(550) xor in_data(549) xor in_data(545) xor in_data(540) xor in_data(539) xor in_data(537) xor in_data(536) xor in_data(535) xor in_data(534) xor in_data(533) xor in_data(532) xor in_data(531) xor in_data(528) xor in_data(527) xor in_data(526) xor in_data(522) xor in_data(521) xor in_data(519) xor in_data(517) xor in_data(514) xor in_data(512) xor in_data(507) xor in_data(502) xor in_data(499) xor in_data(497) xor in_data(496) xor in_data(494) xor in_data(493) xor in_data(492) xor in_data(491) xor in_data(490) xor in_data(488) xor in_data(486) xor in_data(485) xor in_data(484) xor in_data(480) xor in_data(478) xor in_data(477) xor in_data(476) xor in_data(473) xor in_data(468) xor in_data(467) xor in_data(466) xor in_data(465) xor in_data(464) xor in_data(462) xor in_data(461) xor in_data(459) xor in_data(457) xor in_data(455) xor in_data(451) xor in_data(449) xor in_data(448) xor in_data(447) xor in_data(446) xor in_data(444) xor in_data(443) xor in_data(440) xor in_data(439) xor in_data(438) xor in_data(435) xor in_data(434) xor in_data(433) xor in_data(432) xor in_data(431) xor in_data(425) xor in_data(424) xor in_data(423) xor in_data(420) xor in_data(417) xor in_data(415) xor in_data(413) xor in_data(412) xor in_data(409) xor in_data(407) xor in_data(406) xor in_data(405) xor in_data(404) xor in_data(401) xor in_data(399) xor in_data(398) xor in_data(397) xor in_data(391) xor in_data(389) xor in_data(387) xor in_data(386) xor in_data(384) xor in_data(383) xor in_data(380) xor in_data(379) xor in_data(374) xor in_data(373) xor in_data(371) xor in_data(369) xor in_data(368) xor in_data(366) xor in_data(365) xor in_data(364) xor in_data(362) xor in_data(358) xor in_data(356) xor in_data(354) xor in_data(353) xor in_data(352) xor in_data(351) xor in_data(350) xor in_data(349) xor in_data(347) xor in_data(343) xor in_data(342) xor in_data(341) xor in_data(338) xor in_data(337) xor in_data(335) xor in_data(334) xor in_data(333) xor in_data(330) xor in_data(328) xor in_data(324) xor in_data(323) xor in_data(321) xor in_data(314) xor in_data(313) xor in_data(310) xor in_data(307) xor in_data(303) xor in_data(297) xor in_data(294) xor in_data(293) xor in_data(291) xor in_data(290) xor in_data(288) xor in_data(285) xor in_data(284) xor in_data(283) xor in_data(282) xor in_data(279) xor in_data(278) xor in_data(276) xor in_data(274) xor in_data(272) xor in_data(271) xor in_data(266) xor in_data(264) xor in_data(263) xor in_data(262) xor in_data(260) xor in_data(259) xor in_data(257) xor in_data(253) xor in_data(252) xor in_data(247) xor in_data(244) xor in_data(243) xor in_data(242) xor in_data(241) xor in_data(240) xor in_data(239) xor in_data(238) xor in_data(236) xor in_data(235) xor in_data(234) xor in_data(230) xor in_data(229) xor in_data(228) xor in_data(227) xor in_data(220) xor in_data(219) xor in_data(218) xor in_data(216) xor in_data(215) xor in_data(213) xor in_data(212) xor in_data(208) xor in_data(206) xor in_data(202) xor in_data(199) xor in_data(198) xor in_data(195) xor in_data(189) xor in_data(188) xor in_data(186) xor in_data(183) xor in_data(180) xor in_data(179) xor in_data(178) xor in_data(177) xor in_data(175) xor in_data(174) xor in_data(173) xor in_data(172) xor in_data(171) xor in_data(167) xor in_data(165) xor in_data(163) xor in_data(161) xor in_data(160) xor in_data(158) xor in_data(153) xor in_data(151) xor in_data(143) xor in_data(141) xor in_data(140) xor in_data(138) xor in_data(137) xor in_data(135) xor in_data(134) xor in_data(133) xor in_data(132) xor in_data(129) xor in_data(128) xor in_data(127) xor in_data(126) xor in_data(122) xor in_data(118) xor in_data(117) xor in_data(116) xor in_data(115) xor in_data(114) xor in_data(113) xor in_data(111) xor in_data(110) xor in_data(106) xor in_data(105) xor in_data(104) xor in_data(102) xor in_data(100) xor in_data(99) xor in_data(97) xor in_data(95) xor in_data(90) xor in_data(89) xor in_data(86) xor in_data(85) xor in_data(83) xor in_data(82) xor in_data(76) xor in_data(75) xor in_data(66) xor in_data(65) xor in_data(63) xor in_data(62) xor in_data(60) xor in_data(59) xor in_data(57) xor in_data(55) xor in_data(54) xor in_data(53) xor in_data(51) xor in_data(49) xor in_data(48) xor in_data(47) xor in_data(46) xor in_data(41) xor in_data(39) xor in_data(37) xor in_data(34) xor in_data(29) xor in_data(27) xor in_data(26) xor in_data(23) xor in_data(20) xor in_data(19) xor in_data(13) xor in_data(9) xor in_data(6);

out_data(1021)<= in_data(1011) xor in_data(1008) xor in_data(1005) xor in_data(1002) xor in_data(1001) xor in_data(999) xor in_data(996) xor in_data(995) xor in_data(993) xor in_data(991) xor in_data(990) xor in_data(989) xor in_data(988) xor in_data(987) xor in_data(984) xor in_data(983) xor in_data(979) xor in_data(978) xor in_data(977) xor in_data(976) xor in_data(975) xor in_data(972) xor in_data(968) xor in_data(967) xor in_data(966) xor in_data(964) xor in_data(963) xor in_data(962) xor in_data(961) xor in_data(960) xor in_data(959) xor in_data(954) xor in_data(953) xor in_data(952) xor in_data(944) xor in_data(943) xor in_data(942) xor in_data(941) xor in_data(940) xor in_data(939) xor in_data(938) xor in_data(937) xor in_data(936) xor in_data(935) xor in_data(931) xor in_data(930) xor in_data(929) xor in_data(925) xor in_data(922) xor in_data(921) xor in_data(920) xor in_data(918) xor in_data(917) xor in_data(914) xor in_data(912) xor in_data(910) xor in_data(909) xor in_data(908) xor in_data(906) xor in_data(905) xor in_data(904) xor in_data(903) xor in_data(901) xor in_data(899) xor in_data(895) xor in_data(894) xor in_data(893) xor in_data(892) xor in_data(890) xor in_data(887) xor in_data(885) xor in_data(883) xor in_data(877) xor in_data(875) xor in_data(874) xor in_data(873) xor in_data(872) xor in_data(871) xor in_data(870) xor in_data(869) xor in_data(868) xor in_data(866) xor in_data(864) xor in_data(862) xor in_data(860) xor in_data(858) xor in_data(857) xor in_data(856) xor in_data(855) xor in_data(853) xor in_data(848) xor in_data(847) xor in_data(846) xor in_data(844) xor in_data(841) xor in_data(837) xor in_data(836) xor in_data(833) xor in_data(831) xor in_data(830) xor in_data(828) xor in_data(826) xor in_data(825) xor in_data(822) xor in_data(821) xor in_data(820) xor in_data(819) xor in_data(817) xor in_data(815) xor in_data(814) xor in_data(810) xor in_data(809) xor in_data(806) xor in_data(805) xor in_data(804) xor in_data(803) xor in_data(802) xor in_data(801) xor in_data(798) xor in_data(796) xor in_data(794) xor in_data(792) xor in_data(789) xor in_data(788) xor in_data(785) xor in_data(784) xor in_data(781) xor in_data(779) xor in_data(776) xor in_data(775) xor in_data(774) xor in_data(773) xor in_data(772) xor in_data(770) xor in_data(767) xor in_data(766) xor in_data(765) xor in_data(760) xor in_data(756) xor in_data(755) xor in_data(753) xor in_data(752) xor in_data(749) xor in_data(745) xor in_data(743) xor in_data(740) xor in_data(739) xor in_data(737) xor in_data(736) xor in_data(735) xor in_data(734) xor in_data(732) xor in_data(731) xor in_data(730) xor in_data(728) xor in_data(726) xor in_data(724) xor in_data(723) xor in_data(722) xor in_data(719) xor in_data(718) xor in_data(715) xor in_data(714) xor in_data(713) xor in_data(711) xor in_data(710) xor in_data(709) xor in_data(707) xor in_data(706) xor in_data(705) xor in_data(702) xor in_data(701) xor in_data(700) xor in_data(698) xor in_data(696) xor in_data(693) xor in_data(692) xor in_data(691) xor in_data(689) xor in_data(683) xor in_data(682) xor in_data(681) xor in_data(680) xor in_data(678) xor in_data(677) xor in_data(675) xor in_data(674) xor in_data(673) xor in_data(668) xor in_data(667) xor in_data(663) xor in_data(660) xor in_data(658) xor in_data(655) xor in_data(653) xor in_data(652) xor in_data(649) xor in_data(648) xor in_data(646) xor in_data(642) xor in_data(638) xor in_data(636) xor in_data(635) xor in_data(633) xor in_data(630) xor in_data(628) xor in_data(627) xor in_data(626) xor in_data(624) xor in_data(621) xor in_data(620) xor in_data(616) xor in_data(614) xor in_data(613) xor in_data(606) xor in_data(604) xor in_data(601) xor in_data(598) xor in_data(596) xor in_data(595) xor in_data(594) xor in_data(593) xor in_data(592) xor in_data(590) xor in_data(589) xor in_data(588) xor in_data(587) xor in_data(583) xor in_data(582) xor in_data(578) xor in_data(577) xor in_data(575) xor in_data(574) xor in_data(573) xor in_data(571) xor in_data(570) xor in_data(565) xor in_data(564) xor in_data(563) xor in_data(562) xor in_data(559) xor in_data(556) xor in_data(555) xor in_data(554) xor in_data(551) xor in_data(549) xor in_data(548) xor in_data(544) xor in_data(539) xor in_data(538) xor in_data(536) xor in_data(535) xor in_data(534) xor in_data(533) xor in_data(532) xor in_data(531) xor in_data(530) xor in_data(527) xor in_data(526) xor in_data(525) xor in_data(521) xor in_data(520) xor in_data(518) xor in_data(516) xor in_data(513) xor in_data(511) xor in_data(506) xor in_data(501) xor in_data(498) xor in_data(496) xor in_data(495) xor in_data(493) xor in_data(492) xor in_data(491) xor in_data(490) xor in_data(489) xor in_data(487) xor in_data(485) xor in_data(484) xor in_data(483) xor in_data(479) xor in_data(477) xor in_data(476) xor in_data(475) xor in_data(472) xor in_data(467) xor in_data(466) xor in_data(465) xor in_data(464) xor in_data(463) xor in_data(461) xor in_data(460) xor in_data(458) xor in_data(456) xor in_data(454) xor in_data(450) xor in_data(448) xor in_data(447) xor in_data(446) xor in_data(445) xor in_data(443) xor in_data(442) xor in_data(439) xor in_data(438) xor in_data(437) xor in_data(434) xor in_data(433) xor in_data(432) xor in_data(431) xor in_data(430) xor in_data(424) xor in_data(423) xor in_data(422) xor in_data(419) xor in_data(416) xor in_data(414) xor in_data(412) xor in_data(411) xor in_data(408) xor in_data(406) xor in_data(405) xor in_data(404) xor in_data(403) xor in_data(400) xor in_data(398) xor in_data(397) xor in_data(396) xor in_data(390) xor in_data(388) xor in_data(386) xor in_data(385) xor in_data(383) xor in_data(382) xor in_data(379) xor in_data(378) xor in_data(373) xor in_data(372) xor in_data(370) xor in_data(368) xor in_data(367) xor in_data(365) xor in_data(364) xor in_data(363) xor in_data(361) xor in_data(357) xor in_data(355) xor in_data(353) xor in_data(352) xor in_data(351) xor in_data(350) xor in_data(349) xor in_data(348) xor in_data(346) xor in_data(342) xor in_data(341) xor in_data(340) xor in_data(337) xor in_data(336) xor in_data(334) xor in_data(333) xor in_data(332) xor in_data(329) xor in_data(327) xor in_data(323) xor in_data(322) xor in_data(320) xor in_data(313) xor in_data(312) xor in_data(309) xor in_data(306) xor in_data(302) xor in_data(296) xor in_data(293) xor in_data(292) xor in_data(290) xor in_data(289) xor in_data(287) xor in_data(284) xor in_data(283) xor in_data(282) xor in_data(281) xor in_data(278) xor in_data(277) xor in_data(275) xor in_data(273) xor in_data(271) xor in_data(270) xor in_data(265) xor in_data(263) xor in_data(262) xor in_data(261) xor in_data(259) xor in_data(258) xor in_data(256) xor in_data(252) xor in_data(251) xor in_data(246) xor in_data(243) xor in_data(242) xor in_data(241) xor in_data(240) xor in_data(239) xor in_data(238) xor in_data(237) xor in_data(235) xor in_data(234) xor in_data(233) xor in_data(229) xor in_data(228) xor in_data(227) xor in_data(226) xor in_data(219) xor in_data(218) xor in_data(217) xor in_data(215) xor in_data(214) xor in_data(212) xor in_data(211) xor in_data(207) xor in_data(205) xor in_data(201) xor in_data(198) xor in_data(197) xor in_data(194) xor in_data(188) xor in_data(187) xor in_data(185) xor in_data(182) xor in_data(179) xor in_data(178) xor in_data(177) xor in_data(176) xor in_data(174) xor in_data(173) xor in_data(172) xor in_data(171) xor in_data(170) xor in_data(166) xor in_data(164) xor in_data(162) xor in_data(160) xor in_data(159) xor in_data(157) xor in_data(152) xor in_data(150) xor in_data(142) xor in_data(140) xor in_data(139) xor in_data(137) xor in_data(136) xor in_data(134) xor in_data(133) xor in_data(132) xor in_data(131) xor in_data(128) xor in_data(127) xor in_data(126) xor in_data(125) xor in_data(121) xor in_data(117) xor in_data(116) xor in_data(115) xor in_data(114) xor in_data(113) xor in_data(112) xor in_data(110) xor in_data(109) xor in_data(105) xor in_data(104) xor in_data(103) xor in_data(101) xor in_data(99) xor in_data(98) xor in_data(96) xor in_data(94) xor in_data(89) xor in_data(88) xor in_data(85) xor in_data(84) xor in_data(82) xor in_data(81) xor in_data(75) xor in_data(74) xor in_data(65) xor in_data(64) xor in_data(62) xor in_data(61) xor in_data(59) xor in_data(58) xor in_data(56) xor in_data(54) xor in_data(53) xor in_data(52) xor in_data(50) xor in_data(48) xor in_data(47) xor in_data(46) xor in_data(45) xor in_data(40) xor in_data(38) xor in_data(36) xor in_data(33) xor in_data(28) xor in_data(26) xor in_data(25) xor in_data(22) xor in_data(19) xor in_data(18) xor in_data(12) xor in_data(8) xor in_data(5);

out_data(1020)<= in_data(1010) xor in_data(1007) xor in_data(1004) xor in_data(1001) xor in_data(1000) xor in_data(998) xor in_data(995) xor in_data(994) xor in_data(992) xor in_data(990) xor in_data(989) xor in_data(988) xor in_data(987) xor in_data(986) xor in_data(983) xor in_data(982) xor in_data(978) xor in_data(977) xor in_data(976) xor in_data(975) xor in_data(974) xor in_data(971) xor in_data(967) xor in_data(966) xor in_data(965) xor in_data(963) xor in_data(962) xor in_data(961) xor in_data(960) xor in_data(959) xor in_data(958) xor in_data(953) xor in_data(952) xor in_data(951) xor in_data(943) xor in_data(942) xor in_data(941) xor in_data(940) xor in_data(939) xor in_data(938) xor in_data(937) xor in_data(936) xor in_data(935) xor in_data(934) xor in_data(930) xor in_data(929) xor in_data(928) xor in_data(924) xor in_data(921) xor in_data(920) xor in_data(919) xor in_data(917) xor in_data(916) xor in_data(913) xor in_data(911) xor in_data(909) xor in_data(908) xor in_data(907) xor in_data(905) xor in_data(904) xor in_data(903) xor in_data(902) xor in_data(900) xor in_data(898) xor in_data(894) xor in_data(893) xor in_data(892) xor in_data(891) xor in_data(889) xor in_data(886) xor in_data(884) xor in_data(882) xor in_data(876) xor in_data(874) xor in_data(873) xor in_data(872) xor in_data(871) xor in_data(870) xor in_data(869) xor in_data(868) xor in_data(867) xor in_data(865) xor in_data(863) xor in_data(861) xor in_data(859) xor in_data(857) xor in_data(856) xor in_data(855) xor in_data(854) xor in_data(852) xor in_data(847) xor in_data(846) xor in_data(845) xor in_data(843) xor in_data(840) xor in_data(836) xor in_data(835) xor in_data(832) xor in_data(830) xor in_data(829) xor in_data(827) xor in_data(825) xor in_data(824) xor in_data(821) xor in_data(820) xor in_data(819) xor in_data(818) xor in_data(816) xor in_data(814) xor in_data(813) xor in_data(809) xor in_data(808) xor in_data(805) xor in_data(804) xor in_data(803) xor in_data(802) xor in_data(801) xor in_data(800) xor in_data(797) xor in_data(795) xor in_data(793) xor in_data(791) xor in_data(788) xor in_data(787) xor in_data(784) xor in_data(783) xor in_data(780) xor in_data(778) xor in_data(775) xor in_data(774) xor in_data(773) xor in_data(772) xor in_data(771) xor in_data(769) xor in_data(766) xor in_data(765) xor in_data(764) xor in_data(759) xor in_data(755) xor in_data(754) xor in_data(752) xor in_data(751) xor in_data(748) xor in_data(744) xor in_data(742) xor in_data(739) xor in_data(738) xor in_data(736) xor in_data(735) xor in_data(734) xor in_data(733) xor in_data(731) xor in_data(730) xor in_data(729) xor in_data(727) xor in_data(725) xor in_data(723) xor in_data(722) xor in_data(721) xor in_data(718) xor in_data(717) xor in_data(714) xor in_data(713) xor in_data(712) xor in_data(710) xor in_data(709) xor in_data(708) xor in_data(706) xor in_data(705) xor in_data(704) xor in_data(701) xor in_data(700) xor in_data(699) xor in_data(697) xor in_data(695) xor in_data(692) xor in_data(691) xor in_data(690) xor in_data(688) xor in_data(682) xor in_data(681) xor in_data(680) xor in_data(679) xor in_data(677) xor in_data(676) xor in_data(674) xor in_data(673) xor in_data(672) xor in_data(667) xor in_data(666) xor in_data(662) xor in_data(659) xor in_data(657) xor in_data(654) xor in_data(652) xor in_data(651) xor in_data(648) xor in_data(647) xor in_data(645) xor in_data(641) xor in_data(637) xor in_data(635) xor in_data(634) xor in_data(632) xor in_data(629) xor in_data(627) xor in_data(626) xor in_data(625) xor in_data(623) xor in_data(620) xor in_data(619) xor in_data(615) xor in_data(613) xor in_data(612) xor in_data(605) xor in_data(603) xor in_data(600) xor in_data(597) xor in_data(595) xor in_data(594) xor in_data(593) xor in_data(592) xor in_data(591) xor in_data(589) xor in_data(588) xor in_data(587) xor in_data(586) xor in_data(582) xor in_data(581) xor in_data(577) xor in_data(576) xor in_data(574) xor in_data(573) xor in_data(572) xor in_data(570) xor in_data(569) xor in_data(564) xor in_data(563) xor in_data(562) xor in_data(561) xor in_data(558) xor in_data(555) xor in_data(554) xor in_data(553) xor in_data(550) xor in_data(548) xor in_data(547) xor in_data(543) xor in_data(538) xor in_data(537) xor in_data(535) xor in_data(534) xor in_data(533) xor in_data(532) xor in_data(531) xor in_data(530) xor in_data(529) xor in_data(526) xor in_data(525) xor in_data(524) xor in_data(520) xor in_data(519) xor in_data(517) xor in_data(515) xor in_data(512) xor in_data(510) xor in_data(505) xor in_data(500) xor in_data(497) xor in_data(495) xor in_data(494) xor in_data(492) xor in_data(491) xor in_data(490) xor in_data(489) xor in_data(488) xor in_data(486) xor in_data(484) xor in_data(483) xor in_data(482) xor in_data(478) xor in_data(476) xor in_data(475) xor in_data(474) xor in_data(471) xor in_data(466) xor in_data(465) xor in_data(464) xor in_data(463) xor in_data(462) xor in_data(460) xor in_data(459) xor in_data(457) xor in_data(455) xor in_data(453) xor in_data(449) xor in_data(447) xor in_data(446) xor in_data(445) xor in_data(444) xor in_data(442) xor in_data(441) xor in_data(438) xor in_data(437) xor in_data(436) xor in_data(433) xor in_data(432) xor in_data(431) xor in_data(430) xor in_data(429) xor in_data(423) xor in_data(422) xor in_data(421) xor in_data(418) xor in_data(415) xor in_data(413) xor in_data(411) xor in_data(410) xor in_data(407) xor in_data(405) xor in_data(404) xor in_data(403) xor in_data(402) xor in_data(399) xor in_data(397) xor in_data(396) xor in_data(395) xor in_data(389) xor in_data(387) xor in_data(385) xor in_data(384) xor in_data(382) xor in_data(381) xor in_data(378) xor in_data(377) xor in_data(372) xor in_data(371) xor in_data(369) xor in_data(367) xor in_data(366) xor in_data(364) xor in_data(363) xor in_data(362) xor in_data(360) xor in_data(356) xor in_data(354) xor in_data(352) xor in_data(351) xor in_data(350) xor in_data(349) xor in_data(348) xor in_data(347) xor in_data(345) xor in_data(341) xor in_data(340) xor in_data(339) xor in_data(336) xor in_data(335) xor in_data(333) xor in_data(332) xor in_data(331) xor in_data(328) xor in_data(326) xor in_data(322) xor in_data(321) xor in_data(319) xor in_data(312) xor in_data(311) xor in_data(308) xor in_data(305) xor in_data(301) xor in_data(295) xor in_data(292) xor in_data(291) xor in_data(289) xor in_data(288) xor in_data(286) xor in_data(283) xor in_data(282) xor in_data(281) xor in_data(280) xor in_data(277) xor in_data(276) xor in_data(274) xor in_data(272) xor in_data(270) xor in_data(269) xor in_data(264) xor in_data(262) xor in_data(261) xor in_data(260) xor in_data(258) xor in_data(257) xor in_data(255) xor in_data(251) xor in_data(250) xor in_data(245) xor in_data(242) xor in_data(241) xor in_data(240) xor in_data(239) xor in_data(238) xor in_data(237) xor in_data(236) xor in_data(234) xor in_data(233) xor in_data(232) xor in_data(228) xor in_data(227) xor in_data(226) xor in_data(225) xor in_data(218) xor in_data(217) xor in_data(216) xor in_data(214) xor in_data(213) xor in_data(211) xor in_data(210) xor in_data(206) xor in_data(204) xor in_data(200) xor in_data(197) xor in_data(196) xor in_data(193) xor in_data(187) xor in_data(186) xor in_data(184) xor in_data(181) xor in_data(178) xor in_data(177) xor in_data(176) xor in_data(175) xor in_data(173) xor in_data(172) xor in_data(171) xor in_data(170) xor in_data(169) xor in_data(165) xor in_data(163) xor in_data(161) xor in_data(159) xor in_data(158) xor in_data(156) xor in_data(151) xor in_data(149) xor in_data(141) xor in_data(139) xor in_data(138) xor in_data(136) xor in_data(135) xor in_data(133) xor in_data(132) xor in_data(131) xor in_data(130) xor in_data(127) xor in_data(126) xor in_data(125) xor in_data(124) xor in_data(120) xor in_data(116) xor in_data(115) xor in_data(114) xor in_data(113) xor in_data(112) xor in_data(111) xor in_data(109) xor in_data(108) xor in_data(104) xor in_data(103) xor in_data(102) xor in_data(100) xor in_data(98) xor in_data(97) xor in_data(95) xor in_data(93) xor in_data(88) xor in_data(87) xor in_data(84) xor in_data(83) xor in_data(81) xor in_data(80) xor in_data(74) xor in_data(73) xor in_data(64) xor in_data(63) xor in_data(61) xor in_data(60) xor in_data(58) xor in_data(57) xor in_data(55) xor in_data(53) xor in_data(52) xor in_data(51) xor in_data(49) xor in_data(47) xor in_data(46) xor in_data(45) xor in_data(44) xor in_data(39) xor in_data(37) xor in_data(35) xor in_data(32) xor in_data(27) xor in_data(25) xor in_data(24) xor in_data(21) xor in_data(18) xor in_data(17) xor in_data(11) xor in_data(7) xor in_data(4);

out_data(1019)<= in_data(1009) xor in_data(1006) xor in_data(1003) xor in_data(1000) xor in_data(999) xor in_data(997) xor in_data(994) xor in_data(993) xor in_data(991) xor in_data(989) xor in_data(988) xor in_data(987) xor in_data(986) xor in_data(985) xor in_data(982) xor in_data(981) xor in_data(977) xor in_data(976) xor in_data(975) xor in_data(974) xor in_data(973) xor in_data(970) xor in_data(966) xor in_data(965) xor in_data(964) xor in_data(962) xor in_data(961) xor in_data(960) xor in_data(959) xor in_data(958) xor in_data(957) xor in_data(952) xor in_data(951) xor in_data(950) xor in_data(942) xor in_data(941) xor in_data(940) xor in_data(939) xor in_data(938) xor in_data(937) xor in_data(936) xor in_data(935) xor in_data(934) xor in_data(933) xor in_data(929) xor in_data(928) xor in_data(927) xor in_data(923) xor in_data(920) xor in_data(919) xor in_data(918) xor in_data(916) xor in_data(915) xor in_data(912) xor in_data(910) xor in_data(908) xor in_data(907) xor in_data(906) xor in_data(904) xor in_data(903) xor in_data(902) xor in_data(901) xor in_data(899) xor in_data(897) xor in_data(893) xor in_data(892) xor in_data(891) xor in_data(890) xor in_data(888) xor in_data(885) xor in_data(883) xor in_data(881) xor in_data(875) xor in_data(873) xor in_data(872) xor in_data(871) xor in_data(870) xor in_data(869) xor in_data(868) xor in_data(867) xor in_data(866) xor in_data(864) xor in_data(862) xor in_data(860) xor in_data(858) xor in_data(856) xor in_data(855) xor in_data(854) xor in_data(853) xor in_data(851) xor in_data(846) xor in_data(845) xor in_data(844) xor in_data(842) xor in_data(839) xor in_data(835) xor in_data(834) xor in_data(831) xor in_data(829) xor in_data(828) xor in_data(826) xor in_data(824) xor in_data(823) xor in_data(820) xor in_data(819) xor in_data(818) xor in_data(817) xor in_data(815) xor in_data(813) xor in_data(812) xor in_data(808) xor in_data(807) xor in_data(804) xor in_data(803) xor in_data(802) xor in_data(801) xor in_data(800) xor in_data(799) xor in_data(796) xor in_data(794) xor in_data(792) xor in_data(790) xor in_data(787) xor in_data(786) xor in_data(783) xor in_data(782) xor in_data(779) xor in_data(777) xor in_data(774) xor in_data(773) xor in_data(772) xor in_data(771) xor in_data(770) xor in_data(768) xor in_data(765) xor in_data(764) xor in_data(763) xor in_data(758) xor in_data(754) xor in_data(753) xor in_data(751) xor in_data(750) xor in_data(747) xor in_data(743) xor in_data(741) xor in_data(738) xor in_data(737) xor in_data(735) xor in_data(734) xor in_data(733) xor in_data(732) xor in_data(730) xor in_data(729) xor in_data(728) xor in_data(726) xor in_data(724) xor in_data(722) xor in_data(721) xor in_data(720) xor in_data(717) xor in_data(716) xor in_data(713) xor in_data(712) xor in_data(711) xor in_data(709) xor in_data(708) xor in_data(707) xor in_data(705) xor in_data(704) xor in_data(703) xor in_data(700) xor in_data(699) xor in_data(698) xor in_data(696) xor in_data(694) xor in_data(691) xor in_data(690) xor in_data(689) xor in_data(687) xor in_data(681) xor in_data(680) xor in_data(679) xor in_data(678) xor in_data(676) xor in_data(675) xor in_data(673) xor in_data(672) xor in_data(671) xor in_data(666) xor in_data(665) xor in_data(661) xor in_data(658) xor in_data(656) xor in_data(653) xor in_data(651) xor in_data(650) xor in_data(647) xor in_data(646) xor in_data(644) xor in_data(640) xor in_data(636) xor in_data(634) xor in_data(633) xor in_data(631) xor in_data(628) xor in_data(626) xor in_data(625) xor in_data(624) xor in_data(622) xor in_data(619) xor in_data(618) xor in_data(614) xor in_data(612) xor in_data(611) xor in_data(604) xor in_data(602) xor in_data(599) xor in_data(596) xor in_data(594) xor in_data(593) xor in_data(592) xor in_data(591) xor in_data(590) xor in_data(588) xor in_data(587) xor in_data(586) xor in_data(585) xor in_data(581) xor in_data(580) xor in_data(576) xor in_data(575) xor in_data(573) xor in_data(572) xor in_data(571) xor in_data(569) xor in_data(568) xor in_data(563) xor in_data(562) xor in_data(561) xor in_data(560) xor in_data(557) xor in_data(554) xor in_data(553) xor in_data(552) xor in_data(549) xor in_data(547) xor in_data(546) xor in_data(542) xor in_data(537) xor in_data(536) xor in_data(534) xor in_data(533) xor in_data(532) xor in_data(531) xor in_data(530) xor in_data(529) xor in_data(528) xor in_data(525) xor in_data(524) xor in_data(523) xor in_data(519) xor in_data(518) xor in_data(516) xor in_data(514) xor in_data(511) xor in_data(509) xor in_data(504) xor in_data(499) xor in_data(496) xor in_data(494) xor in_data(493) xor in_data(491) xor in_data(490) xor in_data(489) xor in_data(488) xor in_data(487) xor in_data(485) xor in_data(483) xor in_data(482) xor in_data(481) xor in_data(477) xor in_data(475) xor in_data(474) xor in_data(473) xor in_data(470) xor in_data(465) xor in_data(464) xor in_data(463) xor in_data(462) xor in_data(461) xor in_data(459) xor in_data(458) xor in_data(456) xor in_data(454) xor in_data(452) xor in_data(448) xor in_data(446) xor in_data(445) xor in_data(444) xor in_data(443) xor in_data(441) xor in_data(440) xor in_data(437) xor in_data(436) xor in_data(435) xor in_data(432) xor in_data(431) xor in_data(430) xor in_data(429) xor in_data(428) xor in_data(422) xor in_data(421) xor in_data(420) xor in_data(417) xor in_data(414) xor in_data(412) xor in_data(410) xor in_data(409) xor in_data(406) xor in_data(404) xor in_data(403) xor in_data(402) xor in_data(401) xor in_data(398) xor in_data(396) xor in_data(395) xor in_data(394) xor in_data(388) xor in_data(386) xor in_data(384) xor in_data(383) xor in_data(381) xor in_data(380) xor in_data(377) xor in_data(376) xor in_data(371) xor in_data(370) xor in_data(368) xor in_data(366) xor in_data(365) xor in_data(363) xor in_data(362) xor in_data(361) xor in_data(359) xor in_data(355) xor in_data(353) xor in_data(351) xor in_data(350) xor in_data(349) xor in_data(348) xor in_data(347) xor in_data(346) xor in_data(344) xor in_data(340) xor in_data(339) xor in_data(338) xor in_data(335) xor in_data(334) xor in_data(332) xor in_data(331) xor in_data(330) xor in_data(327) xor in_data(325) xor in_data(321) xor in_data(320) xor in_data(318) xor in_data(311) xor in_data(310) xor in_data(307) xor in_data(304) xor in_data(300) xor in_data(294) xor in_data(291) xor in_data(290) xor in_data(288) xor in_data(287) xor in_data(285) xor in_data(282) xor in_data(281) xor in_data(280) xor in_data(279) xor in_data(276) xor in_data(275) xor in_data(273) xor in_data(271) xor in_data(269) xor in_data(268) xor in_data(263) xor in_data(261) xor in_data(260) xor in_data(259) xor in_data(257) xor in_data(256) xor in_data(254) xor in_data(250) xor in_data(249) xor in_data(244) xor in_data(241) xor in_data(240) xor in_data(239) xor in_data(238) xor in_data(237) xor in_data(236) xor in_data(235) xor in_data(233) xor in_data(232) xor in_data(231) xor in_data(227) xor in_data(226) xor in_data(225) xor in_data(224) xor in_data(217) xor in_data(216) xor in_data(215) xor in_data(213) xor in_data(212) xor in_data(210) xor in_data(209) xor in_data(205) xor in_data(203) xor in_data(199) xor in_data(196) xor in_data(195) xor in_data(192) xor in_data(186) xor in_data(185) xor in_data(183) xor in_data(180) xor in_data(177) xor in_data(176) xor in_data(175) xor in_data(174) xor in_data(172) xor in_data(171) xor in_data(170) xor in_data(169) xor in_data(168) xor in_data(164) xor in_data(162) xor in_data(160) xor in_data(158) xor in_data(157) xor in_data(155) xor in_data(150) xor in_data(148) xor in_data(140) xor in_data(138) xor in_data(137) xor in_data(135) xor in_data(134) xor in_data(132) xor in_data(131) xor in_data(130) xor in_data(129) xor in_data(126) xor in_data(125) xor in_data(124) xor in_data(123) xor in_data(119) xor in_data(115) xor in_data(114) xor in_data(113) xor in_data(112) xor in_data(111) xor in_data(110) xor in_data(108) xor in_data(107) xor in_data(103) xor in_data(102) xor in_data(101) xor in_data(99) xor in_data(97) xor in_data(96) xor in_data(94) xor in_data(92) xor in_data(87) xor in_data(86) xor in_data(83) xor in_data(82) xor in_data(80) xor in_data(79) xor in_data(73) xor in_data(72) xor in_data(63) xor in_data(62) xor in_data(60) xor in_data(59) xor in_data(57) xor in_data(56) xor in_data(54) xor in_data(52) xor in_data(51) xor in_data(50) xor in_data(48) xor in_data(46) xor in_data(45) xor in_data(44) xor in_data(43) xor in_data(38) xor in_data(36) xor in_data(34) xor in_data(31) xor in_data(26) xor in_data(24) xor in_data(23) xor in_data(20) xor in_data(17) xor in_data(16) xor in_data(10) xor in_data(6) xor in_data(3);

out_data(1018)<= in_data(1008) xor in_data(1005) xor in_data(1002) xor in_data(999) xor in_data(998) xor in_data(996) xor in_data(993) xor in_data(992) xor in_data(990) xor in_data(988) xor in_data(987) xor in_data(986) xor in_data(985) xor in_data(984) xor in_data(981) xor in_data(980) xor in_data(976) xor in_data(975) xor in_data(974) xor in_data(973) xor in_data(972) xor in_data(969) xor in_data(965) xor in_data(964) xor in_data(963) xor in_data(961) xor in_data(960) xor in_data(959) xor in_data(958) xor in_data(957) xor in_data(956) xor in_data(951) xor in_data(950) xor in_data(949) xor in_data(941) xor in_data(940) xor in_data(939) xor in_data(938) xor in_data(937) xor in_data(936) xor in_data(935) xor in_data(934) xor in_data(933) xor in_data(932) xor in_data(928) xor in_data(927) xor in_data(926) xor in_data(922) xor in_data(919) xor in_data(918) xor in_data(917) xor in_data(915) xor in_data(914) xor in_data(911) xor in_data(909) xor in_data(907) xor in_data(906) xor in_data(905) xor in_data(903) xor in_data(902) xor in_data(901) xor in_data(900) xor in_data(898) xor in_data(896) xor in_data(892) xor in_data(891) xor in_data(890) xor in_data(889) xor in_data(887) xor in_data(884) xor in_data(882) xor in_data(880) xor in_data(874) xor in_data(872) xor in_data(871) xor in_data(870) xor in_data(869) xor in_data(868) xor in_data(867) xor in_data(866) xor in_data(865) xor in_data(863) xor in_data(861) xor in_data(859) xor in_data(857) xor in_data(855) xor in_data(854) xor in_data(853) xor in_data(852) xor in_data(850) xor in_data(845) xor in_data(844) xor in_data(843) xor in_data(841) xor in_data(838) xor in_data(834) xor in_data(833) xor in_data(830) xor in_data(828) xor in_data(827) xor in_data(825) xor in_data(823) xor in_data(822) xor in_data(819) xor in_data(818) xor in_data(817) xor in_data(816) xor in_data(814) xor in_data(812) xor in_data(811) xor in_data(807) xor in_data(806) xor in_data(803) xor in_data(802) xor in_data(801) xor in_data(800) xor in_data(799) xor in_data(798) xor in_data(795) xor in_data(793) xor in_data(791) xor in_data(789) xor in_data(786) xor in_data(785) xor in_data(782) xor in_data(781) xor in_data(778) xor in_data(776) xor in_data(773) xor in_data(772) xor in_data(771) xor in_data(770) xor in_data(769) xor in_data(767) xor in_data(764) xor in_data(763) xor in_data(762) xor in_data(757) xor in_data(753) xor in_data(752) xor in_data(750) xor in_data(749) xor in_data(746) xor in_data(742) xor in_data(740) xor in_data(737) xor in_data(736) xor in_data(734) xor in_data(733) xor in_data(732) xor in_data(731) xor in_data(729) xor in_data(728) xor in_data(727) xor in_data(725) xor in_data(723) xor in_data(721) xor in_data(720) xor in_data(719) xor in_data(716) xor in_data(715) xor in_data(712) xor in_data(711) xor in_data(710) xor in_data(708) xor in_data(707) xor in_data(706) xor in_data(704) xor in_data(703) xor in_data(702) xor in_data(699) xor in_data(698) xor in_data(697) xor in_data(695) xor in_data(693) xor in_data(690) xor in_data(689) xor in_data(688) xor in_data(686) xor in_data(680) xor in_data(679) xor in_data(678) xor in_data(677) xor in_data(675) xor in_data(674) xor in_data(672) xor in_data(671) xor in_data(670) xor in_data(665) xor in_data(664) xor in_data(660) xor in_data(657) xor in_data(655) xor in_data(652) xor in_data(650) xor in_data(649) xor in_data(646) xor in_data(645) xor in_data(643) xor in_data(639) xor in_data(635) xor in_data(633) xor in_data(632) xor in_data(630) xor in_data(627) xor in_data(625) xor in_data(624) xor in_data(623) xor in_data(621) xor in_data(618) xor in_data(617) xor in_data(613) xor in_data(611) xor in_data(610) xor in_data(603) xor in_data(601) xor in_data(598) xor in_data(595) xor in_data(593) xor in_data(592) xor in_data(591) xor in_data(590) xor in_data(589) xor in_data(587) xor in_data(586) xor in_data(585) xor in_data(584) xor in_data(580) xor in_data(579) xor in_data(575) xor in_data(574) xor in_data(572) xor in_data(571) xor in_data(570) xor in_data(568) xor in_data(567) xor in_data(562) xor in_data(561) xor in_data(560) xor in_data(559) xor in_data(556) xor in_data(553) xor in_data(552) xor in_data(551) xor in_data(548) xor in_data(546) xor in_data(545) xor in_data(541) xor in_data(536) xor in_data(535) xor in_data(533) xor in_data(532) xor in_data(531) xor in_data(530) xor in_data(529) xor in_data(528) xor in_data(527) xor in_data(524) xor in_data(523) xor in_data(522) xor in_data(518) xor in_data(517) xor in_data(515) xor in_data(513) xor in_data(510) xor in_data(508) xor in_data(503) xor in_data(498) xor in_data(495) xor in_data(493) xor in_data(492) xor in_data(490) xor in_data(489) xor in_data(488) xor in_data(487) xor in_data(486) xor in_data(484) xor in_data(482) xor in_data(481) xor in_data(480) xor in_data(476) xor in_data(474) xor in_data(473) xor in_data(472) xor in_data(469) xor in_data(464) xor in_data(463) xor in_data(462) xor in_data(461) xor in_data(460) xor in_data(458) xor in_data(457) xor in_data(455) xor in_data(453) xor in_data(451) xor in_data(447) xor in_data(445) xor in_data(444) xor in_data(443) xor in_data(442) xor in_data(440) xor in_data(439) xor in_data(436) xor in_data(435) xor in_data(434) xor in_data(431) xor in_data(430) xor in_data(429) xor in_data(428) xor in_data(427) xor in_data(421) xor in_data(420) xor in_data(419) xor in_data(416) xor in_data(413) xor in_data(411) xor in_data(409) xor in_data(408) xor in_data(405) xor in_data(403) xor in_data(402) xor in_data(401) xor in_data(400) xor in_data(397) xor in_data(395) xor in_data(394) xor in_data(393) xor in_data(387) xor in_data(385) xor in_data(383) xor in_data(382) xor in_data(380) xor in_data(379) xor in_data(376) xor in_data(375) xor in_data(370) xor in_data(369) xor in_data(367) xor in_data(365) xor in_data(364) xor in_data(362) xor in_data(361) xor in_data(360) xor in_data(358) xor in_data(354) xor in_data(352) xor in_data(350) xor in_data(349) xor in_data(348) xor in_data(347) xor in_data(346) xor in_data(345) xor in_data(343) xor in_data(339) xor in_data(338) xor in_data(337) xor in_data(334) xor in_data(333) xor in_data(331) xor in_data(330) xor in_data(329) xor in_data(326) xor in_data(324) xor in_data(320) xor in_data(319) xor in_data(317) xor in_data(310) xor in_data(309) xor in_data(306) xor in_data(303) xor in_data(299) xor in_data(293) xor in_data(290) xor in_data(289) xor in_data(287) xor in_data(286) xor in_data(284) xor in_data(281) xor in_data(280) xor in_data(279) xor in_data(278) xor in_data(275) xor in_data(274) xor in_data(272) xor in_data(270) xor in_data(268) xor in_data(267) xor in_data(262) xor in_data(260) xor in_data(259) xor in_data(258) xor in_data(256) xor in_data(255) xor in_data(253) xor in_data(249) xor in_data(248) xor in_data(243) xor in_data(240) xor in_data(239) xor in_data(238) xor in_data(237) xor in_data(236) xor in_data(235) xor in_data(234) xor in_data(232) xor in_data(231) xor in_data(230) xor in_data(226) xor in_data(225) xor in_data(224) xor in_data(223) xor in_data(216) xor in_data(215) xor in_data(214) xor in_data(212) xor in_data(211) xor in_data(209) xor in_data(208) xor in_data(204) xor in_data(202) xor in_data(198) xor in_data(195) xor in_data(194) xor in_data(191) xor in_data(185) xor in_data(184) xor in_data(182) xor in_data(179) xor in_data(176) xor in_data(175) xor in_data(174) xor in_data(173) xor in_data(171) xor in_data(170) xor in_data(169) xor in_data(168) xor in_data(167) xor in_data(163) xor in_data(161) xor in_data(159) xor in_data(157) xor in_data(156) xor in_data(154) xor in_data(149) xor in_data(147) xor in_data(139) xor in_data(137) xor in_data(136) xor in_data(134) xor in_data(133) xor in_data(131) xor in_data(130) xor in_data(129) xor in_data(128) xor in_data(125) xor in_data(124) xor in_data(123) xor in_data(122) xor in_data(118) xor in_data(114) xor in_data(113) xor in_data(112) xor in_data(111) xor in_data(110) xor in_data(109) xor in_data(107) xor in_data(106) xor in_data(102) xor in_data(101) xor in_data(100) xor in_data(98) xor in_data(96) xor in_data(95) xor in_data(93) xor in_data(91) xor in_data(86) xor in_data(85) xor in_data(82) xor in_data(81) xor in_data(79) xor in_data(78) xor in_data(72) xor in_data(71) xor in_data(62) xor in_data(61) xor in_data(59) xor in_data(58) xor in_data(56) xor in_data(55) xor in_data(53) xor in_data(51) xor in_data(50) xor in_data(49) xor in_data(47) xor in_data(45) xor in_data(44) xor in_data(43) xor in_data(42) xor in_data(37) xor in_data(35) xor in_data(33) xor in_data(30) xor in_data(25) xor in_data(23) xor in_data(22) xor in_data(19) xor in_data(16) xor in_data(15) xor in_data(9) xor in_data(5) xor in_data(2);

out_data(1017)<= in_data(1007) xor in_data(1004) xor in_data(1001) xor in_data(998) xor in_data(997) xor in_data(995) xor in_data(992) xor in_data(991) xor in_data(989) xor in_data(987) xor in_data(986) xor in_data(985) xor in_data(984) xor in_data(983) xor in_data(980) xor in_data(979) xor in_data(975) xor in_data(974) xor in_data(973) xor in_data(972) xor in_data(971) xor in_data(968) xor in_data(964) xor in_data(963) xor in_data(962) xor in_data(960) xor in_data(959) xor in_data(958) xor in_data(957) xor in_data(956) xor in_data(955) xor in_data(950) xor in_data(949) xor in_data(948) xor in_data(940) xor in_data(939) xor in_data(938) xor in_data(937) xor in_data(936) xor in_data(935) xor in_data(934) xor in_data(933) xor in_data(932) xor in_data(931) xor in_data(927) xor in_data(926) xor in_data(925) xor in_data(921) xor in_data(918) xor in_data(917) xor in_data(916) xor in_data(914) xor in_data(913) xor in_data(910) xor in_data(908) xor in_data(906) xor in_data(905) xor in_data(904) xor in_data(902) xor in_data(901) xor in_data(900) xor in_data(899) xor in_data(897) xor in_data(895) xor in_data(891) xor in_data(890) xor in_data(889) xor in_data(888) xor in_data(886) xor in_data(883) xor in_data(881) xor in_data(879) xor in_data(873) xor in_data(871) xor in_data(870) xor in_data(869) xor in_data(868) xor in_data(867) xor in_data(866) xor in_data(865) xor in_data(864) xor in_data(862) xor in_data(860) xor in_data(858) xor in_data(856) xor in_data(854) xor in_data(853) xor in_data(852) xor in_data(851) xor in_data(849) xor in_data(844) xor in_data(843) xor in_data(842) xor in_data(840) xor in_data(837) xor in_data(833) xor in_data(832) xor in_data(829) xor in_data(827) xor in_data(826) xor in_data(824) xor in_data(822) xor in_data(821) xor in_data(818) xor in_data(817) xor in_data(816) xor in_data(815) xor in_data(813) xor in_data(811) xor in_data(810) xor in_data(806) xor in_data(805) xor in_data(802) xor in_data(801) xor in_data(800) xor in_data(799) xor in_data(798) xor in_data(797) xor in_data(794) xor in_data(792) xor in_data(790) xor in_data(788) xor in_data(785) xor in_data(784) xor in_data(781) xor in_data(780) xor in_data(777) xor in_data(775) xor in_data(772) xor in_data(771) xor in_data(770) xor in_data(769) xor in_data(768) xor in_data(766) xor in_data(763) xor in_data(762) xor in_data(761) xor in_data(756) xor in_data(752) xor in_data(751) xor in_data(749) xor in_data(748) xor in_data(745) xor in_data(741) xor in_data(739) xor in_data(736) xor in_data(735) xor in_data(733) xor in_data(732) xor in_data(731) xor in_data(730) xor in_data(728) xor in_data(727) xor in_data(726) xor in_data(724) xor in_data(722) xor in_data(720) xor in_data(719) xor in_data(718) xor in_data(715) xor in_data(714) xor in_data(711) xor in_data(710) xor in_data(709) xor in_data(707) xor in_data(706) xor in_data(705) xor in_data(703) xor in_data(702) xor in_data(701) xor in_data(698) xor in_data(697) xor in_data(696) xor in_data(694) xor in_data(692) xor in_data(689) xor in_data(688) xor in_data(687) xor in_data(685) xor in_data(679) xor in_data(678) xor in_data(677) xor in_data(676) xor in_data(674) xor in_data(673) xor in_data(671) xor in_data(670) xor in_data(669) xor in_data(664) xor in_data(663) xor in_data(659) xor in_data(656) xor in_data(654) xor in_data(651) xor in_data(649) xor in_data(648) xor in_data(645) xor in_data(644) xor in_data(642) xor in_data(638) xor in_data(634) xor in_data(632) xor in_data(631) xor in_data(629) xor in_data(626) xor in_data(624) xor in_data(623) xor in_data(622) xor in_data(620) xor in_data(617) xor in_data(616) xor in_data(612) xor in_data(610) xor in_data(609) xor in_data(602) xor in_data(600) xor in_data(597) xor in_data(594) xor in_data(592) xor in_data(591) xor in_data(590) xor in_data(589) xor in_data(588) xor in_data(586) xor in_data(585) xor in_data(584) xor in_data(583) xor in_data(579) xor in_data(578) xor in_data(574) xor in_data(573) xor in_data(571) xor in_data(570) xor in_data(569) xor in_data(567) xor in_data(566) xor in_data(561) xor in_data(560) xor in_data(559) xor in_data(558) xor in_data(555) xor in_data(552) xor in_data(551) xor in_data(550) xor in_data(547) xor in_data(545) xor in_data(544) xor in_data(540) xor in_data(535) xor in_data(534) xor in_data(532) xor in_data(531) xor in_data(530) xor in_data(529) xor in_data(528) xor in_data(527) xor in_data(526) xor in_data(523) xor in_data(522) xor in_data(521) xor in_data(517) xor in_data(516) xor in_data(514) xor in_data(512) xor in_data(509) xor in_data(507) xor in_data(502) xor in_data(497) xor in_data(494) xor in_data(492) xor in_data(491) xor in_data(489) xor in_data(488) xor in_data(487) xor in_data(486) xor in_data(485) xor in_data(483) xor in_data(481) xor in_data(480) xor in_data(479) xor in_data(475) xor in_data(473) xor in_data(472) xor in_data(471) xor in_data(468) xor in_data(463) xor in_data(462) xor in_data(461) xor in_data(460) xor in_data(459) xor in_data(457) xor in_data(456) xor in_data(454) xor in_data(452) xor in_data(450) xor in_data(446) xor in_data(444) xor in_data(443) xor in_data(442) xor in_data(441) xor in_data(439) xor in_data(438) xor in_data(435) xor in_data(434) xor in_data(433) xor in_data(430) xor in_data(429) xor in_data(428) xor in_data(427) xor in_data(426) xor in_data(420) xor in_data(419) xor in_data(418) xor in_data(415) xor in_data(412) xor in_data(410) xor in_data(408) xor in_data(407) xor in_data(404) xor in_data(402) xor in_data(401) xor in_data(400) xor in_data(399) xor in_data(396) xor in_data(394) xor in_data(393) xor in_data(392) xor in_data(386) xor in_data(384) xor in_data(382) xor in_data(381) xor in_data(379) xor in_data(378) xor in_data(375) xor in_data(374) xor in_data(369) xor in_data(368) xor in_data(366) xor in_data(364) xor in_data(363) xor in_data(361) xor in_data(360) xor in_data(359) xor in_data(357) xor in_data(353) xor in_data(351) xor in_data(349) xor in_data(348) xor in_data(347) xor in_data(346) xor in_data(345) xor in_data(344) xor in_data(342) xor in_data(338) xor in_data(337) xor in_data(336) xor in_data(333) xor in_data(332) xor in_data(330) xor in_data(329) xor in_data(328) xor in_data(325) xor in_data(323) xor in_data(319) xor in_data(318) xor in_data(316) xor in_data(309) xor in_data(308) xor in_data(305) xor in_data(302) xor in_data(298) xor in_data(292) xor in_data(289) xor in_data(288) xor in_data(286) xor in_data(285) xor in_data(283) xor in_data(280) xor in_data(279) xor in_data(278) xor in_data(277) xor in_data(274) xor in_data(273) xor in_data(271) xor in_data(269) xor in_data(267) xor in_data(266) xor in_data(261) xor in_data(259) xor in_data(258) xor in_data(257) xor in_data(255) xor in_data(254) xor in_data(252) xor in_data(248) xor in_data(247) xor in_data(242) xor in_data(239) xor in_data(238) xor in_data(237) xor in_data(236) xor in_data(235) xor in_data(234) xor in_data(233) xor in_data(231) xor in_data(230) xor in_data(229) xor in_data(225) xor in_data(224) xor in_data(223) xor in_data(222) xor in_data(215) xor in_data(214) xor in_data(213) xor in_data(211) xor in_data(210) xor in_data(208) xor in_data(207) xor in_data(203) xor in_data(201) xor in_data(197) xor in_data(194) xor in_data(193) xor in_data(190) xor in_data(184) xor in_data(183) xor in_data(181) xor in_data(178) xor in_data(175) xor in_data(174) xor in_data(173) xor in_data(172) xor in_data(170) xor in_data(169) xor in_data(168) xor in_data(167) xor in_data(166) xor in_data(162) xor in_data(160) xor in_data(158) xor in_data(156) xor in_data(155) xor in_data(153) xor in_data(148) xor in_data(146) xor in_data(138) xor in_data(136) xor in_data(135) xor in_data(133) xor in_data(132) xor in_data(130) xor in_data(129) xor in_data(128) xor in_data(127) xor in_data(124) xor in_data(123) xor in_data(122) xor in_data(121) xor in_data(117) xor in_data(113) xor in_data(112) xor in_data(111) xor in_data(110) xor in_data(109) xor in_data(108) xor in_data(106) xor in_data(105) xor in_data(101) xor in_data(100) xor in_data(99) xor in_data(97) xor in_data(95) xor in_data(94) xor in_data(92) xor in_data(90) xor in_data(85) xor in_data(84) xor in_data(81) xor in_data(80) xor in_data(78) xor in_data(77) xor in_data(71) xor in_data(70) xor in_data(61) xor in_data(60) xor in_data(58) xor in_data(57) xor in_data(55) xor in_data(54) xor in_data(52) xor in_data(50) xor in_data(49) xor in_data(48) xor in_data(46) xor in_data(44) xor in_data(43) xor in_data(42) xor in_data(41) xor in_data(36) xor in_data(34) xor in_data(32) xor in_data(29) xor in_data(24) xor in_data(22) xor in_data(21) xor in_data(18) xor in_data(15) xor in_data(14) xor in_data(8) xor in_data(4) xor in_data(1);

out_data(1016)<= in_data(1006) xor in_data(1003) xor in_data(1000) xor in_data(997) xor in_data(996) xor in_data(994) xor in_data(991) xor in_data(990) xor in_data(988) xor in_data(986) xor in_data(985) xor in_data(984) xor in_data(983) xor in_data(982) xor in_data(979) xor in_data(978) xor in_data(974) xor in_data(973) xor in_data(972) xor in_data(971) xor in_data(970) xor in_data(967) xor in_data(963) xor in_data(962) xor in_data(961) xor in_data(959) xor in_data(958) xor in_data(957) xor in_data(956) xor in_data(955) xor in_data(954) xor in_data(949) xor in_data(948) xor in_data(947) xor in_data(939) xor in_data(938) xor in_data(937) xor in_data(936) xor in_data(935) xor in_data(934) xor in_data(933) xor in_data(932) xor in_data(931) xor in_data(930) xor in_data(926) xor in_data(925) xor in_data(924) xor in_data(920) xor in_data(917) xor in_data(916) xor in_data(915) xor in_data(913) xor in_data(912) xor in_data(909) xor in_data(907) xor in_data(905) xor in_data(904) xor in_data(903) xor in_data(901) xor in_data(900) xor in_data(899) xor in_data(898) xor in_data(896) xor in_data(894) xor in_data(890) xor in_data(889) xor in_data(888) xor in_data(887) xor in_data(885) xor in_data(882) xor in_data(880) xor in_data(878) xor in_data(872) xor in_data(870) xor in_data(869) xor in_data(868) xor in_data(867) xor in_data(866) xor in_data(865) xor in_data(864) xor in_data(863) xor in_data(861) xor in_data(859) xor in_data(857) xor in_data(855) xor in_data(853) xor in_data(852) xor in_data(851) xor in_data(850) xor in_data(848) xor in_data(843) xor in_data(842) xor in_data(841) xor in_data(839) xor in_data(836) xor in_data(832) xor in_data(831) xor in_data(828) xor in_data(826) xor in_data(825) xor in_data(823) xor in_data(821) xor in_data(820) xor in_data(817) xor in_data(816) xor in_data(815) xor in_data(814) xor in_data(812) xor in_data(810) xor in_data(809) xor in_data(805) xor in_data(804) xor in_data(801) xor in_data(800) xor in_data(799) xor in_data(798) xor in_data(797) xor in_data(796) xor in_data(793) xor in_data(791) xor in_data(789) xor in_data(787) xor in_data(784) xor in_data(783) xor in_data(780) xor in_data(779) xor in_data(776) xor in_data(774) xor in_data(771) xor in_data(770) xor in_data(769) xor in_data(768) xor in_data(767) xor in_data(765) xor in_data(762) xor in_data(761) xor in_data(760) xor in_data(755) xor in_data(751) xor in_data(750) xor in_data(748) xor in_data(747) xor in_data(744) xor in_data(740) xor in_data(738) xor in_data(735) xor in_data(734) xor in_data(732) xor in_data(731) xor in_data(730) xor in_data(729) xor in_data(727) xor in_data(726) xor in_data(725) xor in_data(723) xor in_data(721) xor in_data(719) xor in_data(718) xor in_data(717) xor in_data(714) xor in_data(713) xor in_data(710) xor in_data(709) xor in_data(708) xor in_data(706) xor in_data(705) xor in_data(704) xor in_data(702) xor in_data(701) xor in_data(700) xor in_data(697) xor in_data(696) xor in_data(695) xor in_data(693) xor in_data(691) xor in_data(688) xor in_data(687) xor in_data(686) xor in_data(684) xor in_data(678) xor in_data(677) xor in_data(676) xor in_data(675) xor in_data(673) xor in_data(672) xor in_data(670) xor in_data(669) xor in_data(668) xor in_data(663) xor in_data(662) xor in_data(658) xor in_data(655) xor in_data(653) xor in_data(650) xor in_data(648) xor in_data(647) xor in_data(644) xor in_data(643) xor in_data(641) xor in_data(637) xor in_data(633) xor in_data(631) xor in_data(630) xor in_data(628) xor in_data(625) xor in_data(623) xor in_data(622) xor in_data(621) xor in_data(619) xor in_data(616) xor in_data(615) xor in_data(611) xor in_data(609) xor in_data(608) xor in_data(601) xor in_data(599) xor in_data(596) xor in_data(593) xor in_data(591) xor in_data(590) xor in_data(589) xor in_data(588) xor in_data(587) xor in_data(585) xor in_data(584) xor in_data(583) xor in_data(582) xor in_data(578) xor in_data(577) xor in_data(573) xor in_data(572) xor in_data(570) xor in_data(569) xor in_data(568) xor in_data(566) xor in_data(565) xor in_data(560) xor in_data(559) xor in_data(558) xor in_data(557) xor in_data(554) xor in_data(551) xor in_data(550) xor in_data(549) xor in_data(546) xor in_data(544) xor in_data(543) xor in_data(539) xor in_data(534) xor in_data(533) xor in_data(531) xor in_data(530) xor in_data(529) xor in_data(528) xor in_data(527) xor in_data(526) xor in_data(525) xor in_data(522) xor in_data(521) xor in_data(520) xor in_data(516) xor in_data(515) xor in_data(513) xor in_data(511) xor in_data(508) xor in_data(506) xor in_data(501) xor in_data(496) xor in_data(493) xor in_data(491) xor in_data(490) xor in_data(488) xor in_data(487) xor in_data(486) xor in_data(485) xor in_data(484) xor in_data(482) xor in_data(480) xor in_data(479) xor in_data(478) xor in_data(474) xor in_data(472) xor in_data(471) xor in_data(470) xor in_data(467) xor in_data(462) xor in_data(461) xor in_data(460) xor in_data(459) xor in_data(458) xor in_data(456) xor in_data(455) xor in_data(453) xor in_data(451) xor in_data(449) xor in_data(445) xor in_data(443) xor in_data(442) xor in_data(441) xor in_data(440) xor in_data(438) xor in_data(437) xor in_data(434) xor in_data(433) xor in_data(432) xor in_data(429) xor in_data(428) xor in_data(427) xor in_data(426) xor in_data(425) xor in_data(419) xor in_data(418) xor in_data(417) xor in_data(414) xor in_data(411) xor in_data(409) xor in_data(407) xor in_data(406) xor in_data(403) xor in_data(401) xor in_data(400) xor in_data(399) xor in_data(398) xor in_data(395) xor in_data(393) xor in_data(392) xor in_data(391) xor in_data(385) xor in_data(383) xor in_data(381) xor in_data(380) xor in_data(378) xor in_data(377) xor in_data(374) xor in_data(373) xor in_data(368) xor in_data(367) xor in_data(365) xor in_data(363) xor in_data(362) xor in_data(360) xor in_data(359) xor in_data(358) xor in_data(356) xor in_data(352) xor in_data(350) xor in_data(348) xor in_data(347) xor in_data(346) xor in_data(345) xor in_data(344) xor in_data(343) xor in_data(341) xor in_data(337) xor in_data(336) xor in_data(335) xor in_data(332) xor in_data(331) xor in_data(329) xor in_data(328) xor in_data(327) xor in_data(324) xor in_data(322) xor in_data(318) xor in_data(317) xor in_data(315) xor in_data(308) xor in_data(307) xor in_data(304) xor in_data(301) xor in_data(297) xor in_data(291) xor in_data(288) xor in_data(287) xor in_data(285) xor in_data(284) xor in_data(282) xor in_data(279) xor in_data(278) xor in_data(277) xor in_data(276) xor in_data(273) xor in_data(272) xor in_data(270) xor in_data(268) xor in_data(266) xor in_data(265) xor in_data(260) xor in_data(258) xor in_data(257) xor in_data(256) xor in_data(254) xor in_data(253) xor in_data(251) xor in_data(247) xor in_data(246) xor in_data(241) xor in_data(238) xor in_data(237) xor in_data(236) xor in_data(235) xor in_data(234) xor in_data(233) xor in_data(232) xor in_data(230) xor in_data(229) xor in_data(228) xor in_data(224) xor in_data(223) xor in_data(222) xor in_data(221) xor in_data(214) xor in_data(213) xor in_data(212) xor in_data(210) xor in_data(209) xor in_data(207) xor in_data(206) xor in_data(202) xor in_data(200) xor in_data(196) xor in_data(193) xor in_data(192) xor in_data(189) xor in_data(183) xor in_data(182) xor in_data(180) xor in_data(177) xor in_data(174) xor in_data(173) xor in_data(172) xor in_data(171) xor in_data(169) xor in_data(168) xor in_data(167) xor in_data(166) xor in_data(165) xor in_data(161) xor in_data(159) xor in_data(157) xor in_data(155) xor in_data(154) xor in_data(152) xor in_data(147) xor in_data(145) xor in_data(137) xor in_data(135) xor in_data(134) xor in_data(132) xor in_data(131) xor in_data(129) xor in_data(128) xor in_data(127) xor in_data(126) xor in_data(123) xor in_data(122) xor in_data(121) xor in_data(120) xor in_data(116) xor in_data(112) xor in_data(111) xor in_data(110) xor in_data(109) xor in_data(108) xor in_data(107) xor in_data(105) xor in_data(104) xor in_data(100) xor in_data(99) xor in_data(98) xor in_data(96) xor in_data(94) xor in_data(93) xor in_data(91) xor in_data(89) xor in_data(84) xor in_data(83) xor in_data(80) xor in_data(79) xor in_data(77) xor in_data(76) xor in_data(70) xor in_data(69) xor in_data(60) xor in_data(59) xor in_data(57) xor in_data(56) xor in_data(54) xor in_data(53) xor in_data(51) xor in_data(49) xor in_data(48) xor in_data(47) xor in_data(45) xor in_data(43) xor in_data(42) xor in_data(41) xor in_data(40) xor in_data(35) xor in_data(33) xor in_data(31) xor in_data(28) xor in_data(23) xor in_data(21) xor in_data(20) xor in_data(17) xor in_data(14) xor in_data(13) xor in_data(7) xor in_data(3) xor in_data(0);

out_data(1015)<= in_data(1012) xor in_data(1009) xor in_data(1006) xor in_data(1005) xor in_data(1003) xor in_data(1000) xor in_data(999) xor in_data(997) xor in_data(995) xor in_data(994) xor in_data(993) xor in_data(992) xor in_data(991) xor in_data(988) xor in_data(987) xor in_data(983) xor in_data(982) xor in_data(981) xor in_data(980) xor in_data(979) xor in_data(976) xor in_data(972) xor in_data(971) xor in_data(970) xor in_data(968) xor in_data(967) xor in_data(966) xor in_data(965) xor in_data(964) xor in_data(963) xor in_data(958) xor in_data(957) xor in_data(956) xor in_data(948) xor in_data(947) xor in_data(946) xor in_data(945) xor in_data(944) xor in_data(943) xor in_data(942) xor in_data(941) xor in_data(940) xor in_data(939) xor in_data(935) xor in_data(934) xor in_data(933) xor in_data(929) xor in_data(926) xor in_data(925) xor in_data(924) xor in_data(922) xor in_data(921) xor in_data(918) xor in_data(916) xor in_data(914) xor in_data(913) xor in_data(912) xor in_data(910) xor in_data(909) xor in_data(908) xor in_data(907) xor in_data(905) xor in_data(903) xor in_data(899) xor in_data(898) xor in_data(897) xor in_data(896) xor in_data(894) xor in_data(891) xor in_data(889) xor in_data(887) xor in_data(881) xor in_data(879) xor in_data(878) xor in_data(877) xor in_data(876) xor in_data(875) xor in_data(874) xor in_data(873) xor in_data(872) xor in_data(870) xor in_data(868) xor in_data(866) xor in_data(864) xor in_data(862) xor in_data(861) xor in_data(860) xor in_data(859) xor in_data(857) xor in_data(852) xor in_data(851) xor in_data(850) xor in_data(848) xor in_data(845) xor in_data(841) xor in_data(840) xor in_data(837) xor in_data(835) xor in_data(834) xor in_data(832) xor in_data(830) xor in_data(829) xor in_data(826) xor in_data(825) xor in_data(824) xor in_data(823) xor in_data(821) xor in_data(819) xor in_data(818) xor in_data(814) xor in_data(813) xor in_data(810) xor in_data(809) xor in_data(808) xor in_data(807) xor in_data(806) xor in_data(805) xor in_data(802) xor in_data(800) xor in_data(798) xor in_data(796) xor in_data(793) xor in_data(792) xor in_data(789) xor in_data(788) xor in_data(785) xor in_data(783) xor in_data(780) xor in_data(779) xor in_data(778) xor in_data(777) xor in_data(776) xor in_data(774) xor in_data(771) xor in_data(770) xor in_data(769) xor in_data(764) xor in_data(760) xor in_data(759) xor in_data(757) xor in_data(756) xor in_data(753) xor in_data(749) xor in_data(747) xor in_data(744) xor in_data(743) xor in_data(741) xor in_data(740) xor in_data(739) xor in_data(738) xor in_data(736) xor in_data(735) xor in_data(734) xor in_data(732) xor in_data(730) xor in_data(728) xor in_data(727) xor in_data(726) xor in_data(723) xor in_data(722) xor in_data(719) xor in_data(718) xor in_data(717) xor in_data(715) xor in_data(714) xor in_data(713) xor in_data(711) xor in_data(710) xor in_data(709) xor in_data(706) xor in_data(705) xor in_data(704) xor in_data(702) xor in_data(700) xor in_data(697) xor in_data(696) xor in_data(695) xor in_data(693) xor in_data(687) xor in_data(686) xor in_data(685) xor in_data(684) xor in_data(682) xor in_data(681) xor in_data(679) xor in_data(678) xor in_data(677) xor in_data(672) xor in_data(671) xor in_data(667) xor in_data(664) xor in_data(662) xor in_data(659) xor in_data(657) xor in_data(656) xor in_data(653) xor in_data(652) xor in_data(650) xor in_data(646) xor in_data(642) xor in_data(640) xor in_data(639) xor in_data(637) xor in_data(634) xor in_data(632) xor in_data(631) xor in_data(630) xor in_data(628) xor in_data(625) xor in_data(624) xor in_data(620) xor in_data(618) xor in_data(617) xor in_data(610) xor in_data(608) xor in_data(605) xor in_data(602) xor in_data(600) xor in_data(599) xor in_data(598) xor in_data(597) xor in_data(596) xor in_data(594) xor in_data(593) xor in_data(592) xor in_data(591) xor in_data(587) xor in_data(586) xor in_data(582) xor in_data(581) xor in_data(579) xor in_data(578) xor in_data(577) xor in_data(575) xor in_data(574) xor in_data(569) xor in_data(568) xor in_data(567) xor in_data(566) xor in_data(563) xor in_data(560) xor in_data(559) xor in_data(558) xor in_data(555) xor in_data(553) xor in_data(552) xor in_data(548) xor in_data(543) xor in_data(542) xor in_data(540) xor in_data(539) xor in_data(538) xor in_data(537) xor in_data(536) xor in_data(535) xor in_data(534) xor in_data(531) xor in_data(530) xor in_data(529) xor in_data(525) xor in_data(524) xor in_data(522) xor in_data(520) xor in_data(517) xor in_data(515) xor in_data(510) xor in_data(505) xor in_data(502) xor in_data(500) xor in_data(499) xor in_data(497) xor in_data(496) xor in_data(495) xor in_data(494) xor in_data(493) xor in_data(491) xor in_data(489) xor in_data(488) xor in_data(487) xor in_data(483) xor in_data(481) xor in_data(480) xor in_data(479) xor in_data(476) xor in_data(471) xor in_data(470) xor in_data(469) xor in_data(468) xor in_data(467) xor in_data(465) xor in_data(464) xor in_data(462) xor in_data(460) xor in_data(458) xor in_data(454) xor in_data(452) xor in_data(451) xor in_data(450) xor in_data(449) xor in_data(447) xor in_data(446) xor in_data(443) xor in_data(442) xor in_data(441) xor in_data(438) xor in_data(437) xor in_data(436) xor in_data(435) xor in_data(434) xor in_data(428) xor in_data(427) xor in_data(426) xor in_data(423) xor in_data(420) xor in_data(418) xor in_data(416) xor in_data(415) xor in_data(412) xor in_data(410) xor in_data(409) xor in_data(408) xor in_data(407) xor in_data(404) xor in_data(402) xor in_data(401) xor in_data(400) xor in_data(394) xor in_data(392) xor in_data(390) xor in_data(389) xor in_data(387) xor in_data(386) xor in_data(383) xor in_data(382) xor in_data(377) xor in_data(376) xor in_data(374) xor in_data(372) xor in_data(371) xor in_data(369) xor in_data(368) xor in_data(367) xor in_data(365) xor in_data(361) xor in_data(359) xor in_data(357) xor in_data(356) xor in_data(355) xor in_data(354) xor in_data(353) xor in_data(352) xor in_data(350) xor in_data(346) xor in_data(345) xor in_data(344) xor in_data(341) xor in_data(340) xor in_data(338) xor in_data(337) xor in_data(336) xor in_data(333) xor in_data(331) xor in_data(327) xor in_data(326) xor in_data(324) xor in_data(317) xor in_data(316) xor in_data(313) xor in_data(310) xor in_data(306) xor in_data(300) xor in_data(297) xor in_data(296) xor in_data(294) xor in_data(293) xor in_data(291) xor in_data(288) xor in_data(287) xor in_data(286) xor in_data(285) xor in_data(282) xor in_data(281) xor in_data(279) xor in_data(277) xor in_data(275) xor in_data(274) xor in_data(269) xor in_data(267) xor in_data(266) xor in_data(265) xor in_data(263) xor in_data(262) xor in_data(260) xor in_data(256) xor in_data(255) xor in_data(250) xor in_data(247) xor in_data(246) xor in_data(245) xor in_data(244) xor in_data(243) xor in_data(242) xor in_data(241) xor in_data(239) xor in_data(238) xor in_data(237) xor in_data(233) xor in_data(232) xor in_data(231) xor in_data(230) xor in_data(223) xor in_data(222) xor in_data(221) xor in_data(219) xor in_data(218) xor in_data(216) xor in_data(215) xor in_data(211) xor in_data(209) xor in_data(205) xor in_data(202) xor in_data(201) xor in_data(198) xor in_data(192) xor in_data(191) xor in_data(189) xor in_data(186) xor in_data(183) xor in_data(182) xor in_data(181) xor in_data(180) xor in_data(178) xor in_data(177) xor in_data(176) xor in_data(175) xor in_data(174) xor in_data(170) xor in_data(168) xor in_data(166) xor in_data(164) xor in_data(163) xor in_data(161) xor in_data(156) xor in_data(154) xor in_data(146) xor in_data(144) xor in_data(143) xor in_data(141) xor in_data(140) xor in_data(138) xor in_data(137) xor in_data(136) xor in_data(135) xor in_data(132) xor in_data(131) xor in_data(130) xor in_data(129) xor in_data(125) xor in_data(121) xor in_data(120) xor in_data(119) xor in_data(118) xor in_data(117) xor in_data(116) xor in_data(114) xor in_data(113) xor in_data(109) xor in_data(108) xor in_data(107) xor in_data(105) xor in_data(103) xor in_data(102) xor in_data(100) xor in_data(98) xor in_data(93) xor in_data(92) xor in_data(89) xor in_data(88) xor in_data(86) xor in_data(85) xor in_data(79) xor in_data(78) xor in_data(69) xor in_data(68) xor in_data(66) xor in_data(65) xor in_data(63) xor in_data(62) xor in_data(60) xor in_data(58) xor in_data(57) xor in_data(56) xor in_data(54) xor in_data(52) xor in_data(51) xor in_data(50) xor in_data(49) xor in_data(44) xor in_data(42) xor in_data(40) xor in_data(37) xor in_data(32) xor in_data(30) xor in_data(29) xor in_data(26) xor in_data(23) xor in_data(22) xor in_data(16) xor in_data(12) xor in_data(9) xor in_data(2);

out_data(1014)<= in_data(1011) xor in_data(1008) xor in_data(1005) xor in_data(1004) xor in_data(1002) xor in_data(999) xor in_data(998) xor in_data(996) xor in_data(994) xor in_data(993) xor in_data(992) xor in_data(991) xor in_data(990) xor in_data(987) xor in_data(986) xor in_data(982) xor in_data(981) xor in_data(980) xor in_data(979) xor in_data(978) xor in_data(975) xor in_data(971) xor in_data(970) xor in_data(969) xor in_data(967) xor in_data(966) xor in_data(965) xor in_data(964) xor in_data(963) xor in_data(962) xor in_data(957) xor in_data(956) xor in_data(955) xor in_data(947) xor in_data(946) xor in_data(945) xor in_data(944) xor in_data(943) xor in_data(942) xor in_data(941) xor in_data(940) xor in_data(939) xor in_data(938) xor in_data(934) xor in_data(933) xor in_data(932) xor in_data(928) xor in_data(925) xor in_data(924) xor in_data(923) xor in_data(921) xor in_data(920) xor in_data(917) xor in_data(915) xor in_data(913) xor in_data(912) xor in_data(911) xor in_data(909) xor in_data(908) xor in_data(907) xor in_data(906) xor in_data(904) xor in_data(902) xor in_data(898) xor in_data(897) xor in_data(896) xor in_data(895) xor in_data(893) xor in_data(890) xor in_data(888) xor in_data(886) xor in_data(880) xor in_data(878) xor in_data(877) xor in_data(876) xor in_data(875) xor in_data(874) xor in_data(873) xor in_data(872) xor in_data(871) xor in_data(869) xor in_data(867) xor in_data(865) xor in_data(863) xor in_data(861) xor in_data(860) xor in_data(859) xor in_data(858) xor in_data(856) xor in_data(851) xor in_data(850) xor in_data(849) xor in_data(847) xor in_data(844) xor in_data(840) xor in_data(839) xor in_data(836) xor in_data(834) xor in_data(833) xor in_data(831) xor in_data(829) xor in_data(828) xor in_data(825) xor in_data(824) xor in_data(823) xor in_data(822) xor in_data(820) xor in_data(818) xor in_data(817) xor in_data(813) xor in_data(812) xor in_data(809) xor in_data(808) xor in_data(807) xor in_data(806) xor in_data(805) xor in_data(804) xor in_data(801) xor in_data(799) xor in_data(797) xor in_data(795) xor in_data(792) xor in_data(791) xor in_data(788) xor in_data(787) xor in_data(784) xor in_data(782) xor in_data(779) xor in_data(778) xor in_data(777) xor in_data(776) xor in_data(775) xor in_data(773) xor in_data(770) xor in_data(769) xor in_data(768) xor in_data(763) xor in_data(759) xor in_data(758) xor in_data(756) xor in_data(755) xor in_data(752) xor in_data(748) xor in_data(746) xor in_data(743) xor in_data(742) xor in_data(740) xor in_data(739) xor in_data(738) xor in_data(737) xor in_data(735) xor in_data(734) xor in_data(733) xor in_data(731) xor in_data(729) xor in_data(727) xor in_data(726) xor in_data(725) xor in_data(722) xor in_data(721) xor in_data(718) xor in_data(717) xor in_data(716) xor in_data(714) xor in_data(713) xor in_data(712) xor in_data(710) xor in_data(709) xor in_data(708) xor in_data(705) xor in_data(704) xor in_data(703) xor in_data(701) xor in_data(699) xor in_data(696) xor in_data(695) xor in_data(694) xor in_data(692) xor in_data(686) xor in_data(685) xor in_data(684) xor in_data(683) xor in_data(681) xor in_data(680) xor in_data(678) xor in_data(677) xor in_data(676) xor in_data(671) xor in_data(670) xor in_data(666) xor in_data(663) xor in_data(661) xor in_data(658) xor in_data(656) xor in_data(655) xor in_data(652) xor in_data(651) xor in_data(649) xor in_data(645) xor in_data(641) xor in_data(639) xor in_data(638) xor in_data(636) xor in_data(633) xor in_data(631) xor in_data(630) xor in_data(629) xor in_data(627) xor in_data(624) xor in_data(623) xor in_data(619) xor in_data(617) xor in_data(616) xor in_data(609) xor in_data(607) xor in_data(604) xor in_data(601) xor in_data(599) xor in_data(598) xor in_data(597) xor in_data(596) xor in_data(595) xor in_data(593) xor in_data(592) xor in_data(591) xor in_data(590) xor in_data(586) xor in_data(585) xor in_data(581) xor in_data(580) xor in_data(578) xor in_data(577) xor in_data(576) xor in_data(574) xor in_data(573) xor in_data(568) xor in_data(567) xor in_data(566) xor in_data(565) xor in_data(562) xor in_data(559) xor in_data(558) xor in_data(557) xor in_data(554) xor in_data(552) xor in_data(551) xor in_data(547) xor in_data(542) xor in_data(541) xor in_data(539) xor in_data(538) xor in_data(537) xor in_data(536) xor in_data(535) xor in_data(534) xor in_data(533) xor in_data(530) xor in_data(529) xor in_data(528) xor in_data(524) xor in_data(523) xor in_data(521) xor in_data(519) xor in_data(516) xor in_data(514) xor in_data(509) xor in_data(504) xor in_data(501) xor in_data(499) xor in_data(498) xor in_data(496) xor in_data(495) xor in_data(494) xor in_data(493) xor in_data(492) xor in_data(490) xor in_data(488) xor in_data(487) xor in_data(486) xor in_data(482) xor in_data(480) xor in_data(479) xor in_data(478) xor in_data(475) xor in_data(470) xor in_data(469) xor in_data(468) xor in_data(467) xor in_data(466) xor in_data(464) xor in_data(463) xor in_data(461) xor in_data(459) xor in_data(457) xor in_data(453) xor in_data(451) xor in_data(450) xor in_data(449) xor in_data(448) xor in_data(446) xor in_data(445) xor in_data(442) xor in_data(441) xor in_data(440) xor in_data(437) xor in_data(436) xor in_data(435) xor in_data(434) xor in_data(433) xor in_data(427) xor in_data(426) xor in_data(425) xor in_data(422) xor in_data(419) xor in_data(417) xor in_data(415) xor in_data(414) xor in_data(411) xor in_data(409) xor in_data(408) xor in_data(407) xor in_data(406) xor in_data(403) xor in_data(401) xor in_data(400) xor in_data(399) xor in_data(393) xor in_data(391) xor in_data(389) xor in_data(388) xor in_data(386) xor in_data(385) xor in_data(382) xor in_data(381) xor in_data(376) xor in_data(375) xor in_data(373) xor in_data(371) xor in_data(370) xor in_data(368) xor in_data(367) xor in_data(366) xor in_data(364) xor in_data(360) xor in_data(358) xor in_data(356) xor in_data(355) xor in_data(354) xor in_data(353) xor in_data(352) xor in_data(351) xor in_data(349) xor in_data(345) xor in_data(344) xor in_data(343) xor in_data(340) xor in_data(339) xor in_data(337) xor in_data(336) xor in_data(335) xor in_data(332) xor in_data(330) xor in_data(326) xor in_data(325) xor in_data(323) xor in_data(316) xor in_data(315) xor in_data(312) xor in_data(309) xor in_data(305) xor in_data(299) xor in_data(296) xor in_data(295) xor in_data(293) xor in_data(292) xor in_data(290) xor in_data(287) xor in_data(286) xor in_data(285) xor in_data(284) xor in_data(281) xor in_data(280) xor in_data(278) xor in_data(276) xor in_data(274) xor in_data(273) xor in_data(268) xor in_data(266) xor in_data(265) xor in_data(264) xor in_data(262) xor in_data(261) xor in_data(259) xor in_data(255) xor in_data(254) xor in_data(249) xor in_data(246) xor in_data(245) xor in_data(244) xor in_data(243) xor in_data(242) xor in_data(241) xor in_data(240) xor in_data(238) xor in_data(237) xor in_data(236) xor in_data(232) xor in_data(231) xor in_data(230) xor in_data(229) xor in_data(222) xor in_data(221) xor in_data(220) xor in_data(218) xor in_data(217) xor in_data(215) xor in_data(214) xor in_data(210) xor in_data(208) xor in_data(204) xor in_data(201) xor in_data(200) xor in_data(197) xor in_data(191) xor in_data(190) xor in_data(188) xor in_data(185) xor in_data(182) xor in_data(181) xor in_data(180) xor in_data(179) xor in_data(177) xor in_data(176) xor in_data(175) xor in_data(174) xor in_data(173) xor in_data(169) xor in_data(167) xor in_data(165) xor in_data(163) xor in_data(162) xor in_data(160) xor in_data(155) xor in_data(153) xor in_data(145) xor in_data(143) xor in_data(142) xor in_data(140) xor in_data(139) xor in_data(137) xor in_data(136) xor in_data(135) xor in_data(134) xor in_data(131) xor in_data(130) xor in_data(129) xor in_data(128) xor in_data(124) xor in_data(120) xor in_data(119) xor in_data(118) xor in_data(117) xor in_data(116) xor in_data(115) xor in_data(113) xor in_data(112) xor in_data(108) xor in_data(107) xor in_data(106) xor in_data(104) xor in_data(102) xor in_data(101) xor in_data(99) xor in_data(97) xor in_data(92) xor in_data(91) xor in_data(88) xor in_data(87) xor in_data(85) xor in_data(84) xor in_data(78) xor in_data(77) xor in_data(68) xor in_data(67) xor in_data(65) xor in_data(64) xor in_data(62) xor in_data(61) xor in_data(59) xor in_data(57) xor in_data(56) xor in_data(55) xor in_data(53) xor in_data(51) xor in_data(50) xor in_data(49) xor in_data(48) xor in_data(43) xor in_data(41) xor in_data(39) xor in_data(36) xor in_data(31) xor in_data(29) xor in_data(28) xor in_data(25) xor in_data(22) xor in_data(21) xor in_data(15) xor in_data(11) xor in_data(8) xor in_data(1);

out_data(1013)<= in_data(1010) xor in_data(1007) xor in_data(1004) xor in_data(1003) xor in_data(1001) xor in_data(998) xor in_data(997) xor in_data(995) xor in_data(993) xor in_data(992) xor in_data(991) xor in_data(990) xor in_data(989) xor in_data(986) xor in_data(985) xor in_data(981) xor in_data(980) xor in_data(979) xor in_data(978) xor in_data(977) xor in_data(974) xor in_data(970) xor in_data(969) xor in_data(968) xor in_data(966) xor in_data(965) xor in_data(964) xor in_data(963) xor in_data(962) xor in_data(961) xor in_data(956) xor in_data(955) xor in_data(954) xor in_data(946) xor in_data(945) xor in_data(944) xor in_data(943) xor in_data(942) xor in_data(941) xor in_data(940) xor in_data(939) xor in_data(938) xor in_data(937) xor in_data(933) xor in_data(932) xor in_data(931) xor in_data(927) xor in_data(924) xor in_data(923) xor in_data(922) xor in_data(920) xor in_data(919) xor in_data(916) xor in_data(914) xor in_data(912) xor in_data(911) xor in_data(910) xor in_data(908) xor in_data(907) xor in_data(906) xor in_data(905) xor in_data(903) xor in_data(901) xor in_data(897) xor in_data(896) xor in_data(895) xor in_data(894) xor in_data(892) xor in_data(889) xor in_data(887) xor in_data(885) xor in_data(879) xor in_data(877) xor in_data(876) xor in_data(875) xor in_data(874) xor in_data(873) xor in_data(872) xor in_data(871) xor in_data(870) xor in_data(868) xor in_data(866) xor in_data(864) xor in_data(862) xor in_data(860) xor in_data(859) xor in_data(858) xor in_data(857) xor in_data(855) xor in_data(850) xor in_data(849) xor in_data(848) xor in_data(846) xor in_data(843) xor in_data(839) xor in_data(838) xor in_data(835) xor in_data(833) xor in_data(832) xor in_data(830) xor in_data(828) xor in_data(827) xor in_data(824) xor in_data(823) xor in_data(822) xor in_data(821) xor in_data(819) xor in_data(817) xor in_data(816) xor in_data(812) xor in_data(811) xor in_data(808) xor in_data(807) xor in_data(806) xor in_data(805) xor in_data(804) xor in_data(803) xor in_data(800) xor in_data(798) xor in_data(796) xor in_data(794) xor in_data(791) xor in_data(790) xor in_data(787) xor in_data(786) xor in_data(783) xor in_data(781) xor in_data(778) xor in_data(777) xor in_data(776) xor in_data(775) xor in_data(774) xor in_data(772) xor in_data(769) xor in_data(768) xor in_data(767) xor in_data(762) xor in_data(758) xor in_data(757) xor in_data(755) xor in_data(754) xor in_data(751) xor in_data(747) xor in_data(745) xor in_data(742) xor in_data(741) xor in_data(739) xor in_data(738) xor in_data(737) xor in_data(736) xor in_data(734) xor in_data(733) xor in_data(732) xor in_data(730) xor in_data(728) xor in_data(726) xor in_data(725) xor in_data(724) xor in_data(721) xor in_data(720) xor in_data(717) xor in_data(716) xor in_data(715) xor in_data(713) xor in_data(712) xor in_data(711) xor in_data(709) xor in_data(708) xor in_data(707) xor in_data(704) xor in_data(703) xor in_data(702) xor in_data(700) xor in_data(698) xor in_data(695) xor in_data(694) xor in_data(693) xor in_data(691) xor in_data(685) xor in_data(684) xor in_data(683) xor in_data(682) xor in_data(680) xor in_data(679) xor in_data(677) xor in_data(676) xor in_data(675) xor in_data(670) xor in_data(669) xor in_data(665) xor in_data(662) xor in_data(660) xor in_data(657) xor in_data(655) xor in_data(654) xor in_data(651) xor in_data(650) xor in_data(648) xor in_data(644) xor in_data(640) xor in_data(638) xor in_data(637) xor in_data(635) xor in_data(632) xor in_data(630) xor in_data(629) xor in_data(628) xor in_data(626) xor in_data(623) xor in_data(622) xor in_data(618) xor in_data(616) xor in_data(615) xor in_data(608) xor in_data(606) xor in_data(603) xor in_data(600) xor in_data(598) xor in_data(597) xor in_data(596) xor in_data(595) xor in_data(594) xor in_data(592) xor in_data(591) xor in_data(590) xor in_data(589) xor in_data(585) xor in_data(584) xor in_data(580) xor in_data(579) xor in_data(577) xor in_data(576) xor in_data(575) xor in_data(573) xor in_data(572) xor in_data(567) xor in_data(566) xor in_data(565) xor in_data(564) xor in_data(561) xor in_data(558) xor in_data(557) xor in_data(556) xor in_data(553) xor in_data(551) xor in_data(550) xor in_data(546) xor in_data(541) xor in_data(540) xor in_data(538) xor in_data(537) xor in_data(536) xor in_data(535) xor in_data(534) xor in_data(533) xor in_data(532) xor in_data(529) xor in_data(528) xor in_data(527) xor in_data(523) xor in_data(522) xor in_data(520) xor in_data(518) xor in_data(515) xor in_data(513) xor in_data(508) xor in_data(503) xor in_data(500) xor in_data(498) xor in_data(497) xor in_data(495) xor in_data(494) xor in_data(493) xor in_data(492) xor in_data(491) xor in_data(489) xor in_data(487) xor in_data(486) xor in_data(485) xor in_data(481) xor in_data(479) xor in_data(478) xor in_data(477) xor in_data(474) xor in_data(469) xor in_data(468) xor in_data(467) xor in_data(466) xor in_data(465) xor in_data(463) xor in_data(462) xor in_data(460) xor in_data(458) xor in_data(456) xor in_data(452) xor in_data(450) xor in_data(449) xor in_data(448) xor in_data(447) xor in_data(445) xor in_data(444) xor in_data(441) xor in_data(440) xor in_data(439) xor in_data(436) xor in_data(435) xor in_data(434) xor in_data(433) xor in_data(432) xor in_data(426) xor in_data(425) xor in_data(424) xor in_data(421) xor in_data(418) xor in_data(416) xor in_data(414) xor in_data(413) xor in_data(410) xor in_data(408) xor in_data(407) xor in_data(406) xor in_data(405) xor in_data(402) xor in_data(400) xor in_data(399) xor in_data(398) xor in_data(392) xor in_data(390) xor in_data(388) xor in_data(387) xor in_data(385) xor in_data(384) xor in_data(381) xor in_data(380) xor in_data(375) xor in_data(374) xor in_data(372) xor in_data(370) xor in_data(369) xor in_data(367) xor in_data(366) xor in_data(365) xor in_data(363) xor in_data(359) xor in_data(357) xor in_data(355) xor in_data(354) xor in_data(353) xor in_data(352) xor in_data(351) xor in_data(350) xor in_data(348) xor in_data(344) xor in_data(343) xor in_data(342) xor in_data(339) xor in_data(338) xor in_data(336) xor in_data(335) xor in_data(334) xor in_data(331) xor in_data(329) xor in_data(325) xor in_data(324) xor in_data(322) xor in_data(315) xor in_data(314) xor in_data(311) xor in_data(308) xor in_data(304) xor in_data(298) xor in_data(295) xor in_data(294) xor in_data(292) xor in_data(291) xor in_data(289) xor in_data(286) xor in_data(285) xor in_data(284) xor in_data(283) xor in_data(280) xor in_data(279) xor in_data(277) xor in_data(275) xor in_data(273) xor in_data(272) xor in_data(267) xor in_data(265) xor in_data(264) xor in_data(263) xor in_data(261) xor in_data(260) xor in_data(258) xor in_data(254) xor in_data(253) xor in_data(248) xor in_data(245) xor in_data(244) xor in_data(243) xor in_data(242) xor in_data(241) xor in_data(240) xor in_data(239) xor in_data(237) xor in_data(236) xor in_data(235) xor in_data(231) xor in_data(230) xor in_data(229) xor in_data(228) xor in_data(221) xor in_data(220) xor in_data(219) xor in_data(217) xor in_data(216) xor in_data(214) xor in_data(213) xor in_data(209) xor in_data(207) xor in_data(203) xor in_data(200) xor in_data(199) xor in_data(196) xor in_data(190) xor in_data(189) xor in_data(187) xor in_data(184) xor in_data(181) xor in_data(180) xor in_data(179) xor in_data(178) xor in_data(176) xor in_data(175) xor in_data(174) xor in_data(173) xor in_data(172) xor in_data(168) xor in_data(166) xor in_data(164) xor in_data(162) xor in_data(161) xor in_data(159) xor in_data(154) xor in_data(152) xor in_data(144) xor in_data(142) xor in_data(141) xor in_data(139) xor in_data(138) xor in_data(136) xor in_data(135) xor in_data(134) xor in_data(133) xor in_data(130) xor in_data(129) xor in_data(128) xor in_data(127) xor in_data(123) xor in_data(119) xor in_data(118) xor in_data(117) xor in_data(116) xor in_data(115) xor in_data(114) xor in_data(112) xor in_data(111) xor in_data(107) xor in_data(106) xor in_data(105) xor in_data(103) xor in_data(101) xor in_data(100) xor in_data(98) xor in_data(96) xor in_data(91) xor in_data(90) xor in_data(87) xor in_data(86) xor in_data(84) xor in_data(83) xor in_data(77) xor in_data(76) xor in_data(67) xor in_data(66) xor in_data(64) xor in_data(63) xor in_data(61) xor in_data(60) xor in_data(58) xor in_data(56) xor in_data(55) xor in_data(54) xor in_data(52) xor in_data(50) xor in_data(49) xor in_data(48) xor in_data(47) xor in_data(42) xor in_data(40) xor in_data(38) xor in_data(35) xor in_data(30) xor in_data(28) xor in_data(27) xor in_data(24) xor in_data(21) xor in_data(20) xor in_data(14) xor in_data(10) xor in_data(7) xor in_data(0);

end;