library ieee;
use ieee.std_logic_1164.all;
entity chien is
    port(
        a_1     :    in  std_logic_vector(8 downto 0);
        a_2     :    in  std_logic_vector(8 downto 0);
        E     :    out std_logic_vector(510 downto 0)
);
end entity;

architecture arch of chien is
    signal mulr_1_1 : std_logic_vector(8 downto 0);
    signal mulr_2_1 : std_logic_vector(8 downto 0);
    signal mulr_1_2 : std_logic_vector(8 downto 0);
    signal mulr_2_2 : std_logic_vector(8 downto 0);
    signal mulr_1_3 : std_logic_vector(8 downto 0);
    signal mulr_2_3 : std_logic_vector(8 downto 0);
    signal mulr_1_4 : std_logic_vector(8 downto 0);
    signal mulr_2_4 : std_logic_vector(8 downto 0);
    signal mulr_1_5 : std_logic_vector(8 downto 0);
    signal mulr_2_5 : std_logic_vector(8 downto 0);
    signal mulr_1_6 : std_logic_vector(8 downto 0);
    signal mulr_2_6 : std_logic_vector(8 downto 0);
    signal mulr_1_7 : std_logic_vector(8 downto 0);
    signal mulr_2_7 : std_logic_vector(8 downto 0);
    signal mulr_1_8 : std_logic_vector(8 downto 0);
    signal mulr_2_8 : std_logic_vector(8 downto 0);
    signal mulr_1_9 : std_logic_vector(8 downto 0);
    signal mulr_2_9 : std_logic_vector(8 downto 0);
    signal mulr_1_10 : std_logic_vector(8 downto 0);
    signal mulr_2_10 : std_logic_vector(8 downto 0);
    signal mulr_1_11 : std_logic_vector(8 downto 0);
    signal mulr_2_11 : std_logic_vector(8 downto 0);
    signal mulr_1_12 : std_logic_vector(8 downto 0);
    signal mulr_2_12 : std_logic_vector(8 downto 0);
    signal mulr_1_13 : std_logic_vector(8 downto 0);
    signal mulr_2_13 : std_logic_vector(8 downto 0);
    signal mulr_1_14 : std_logic_vector(8 downto 0);
    signal mulr_2_14 : std_logic_vector(8 downto 0);
    signal mulr_1_15 : std_logic_vector(8 downto 0);
    signal mulr_2_15 : std_logic_vector(8 downto 0);
    signal mulr_1_16 : std_logic_vector(8 downto 0);
    signal mulr_2_16 : std_logic_vector(8 downto 0);
    signal mulr_1_17 : std_logic_vector(8 downto 0);
    signal mulr_2_17 : std_logic_vector(8 downto 0);
    signal mulr_1_18 : std_logic_vector(8 downto 0);
    signal mulr_2_18 : std_logic_vector(8 downto 0);
    signal mulr_1_19 : std_logic_vector(8 downto 0);
    signal mulr_2_19 : std_logic_vector(8 downto 0);
    signal mulr_1_20 : std_logic_vector(8 downto 0);
    signal mulr_2_20 : std_logic_vector(8 downto 0);
    signal mulr_1_21 : std_logic_vector(8 downto 0);
    signal mulr_2_21 : std_logic_vector(8 downto 0);
    signal mulr_1_22 : std_logic_vector(8 downto 0);
    signal mulr_2_22 : std_logic_vector(8 downto 0);
    signal mulr_1_23 : std_logic_vector(8 downto 0);
    signal mulr_2_23 : std_logic_vector(8 downto 0);
    signal mulr_1_24 : std_logic_vector(8 downto 0);
    signal mulr_2_24 : std_logic_vector(8 downto 0);
    signal mulr_1_25 : std_logic_vector(8 downto 0);
    signal mulr_2_25 : std_logic_vector(8 downto 0);
    signal mulr_1_26 : std_logic_vector(8 downto 0);
    signal mulr_2_26 : std_logic_vector(8 downto 0);
    signal mulr_1_27 : std_logic_vector(8 downto 0);
    signal mulr_2_27 : std_logic_vector(8 downto 0);
    signal mulr_1_28 : std_logic_vector(8 downto 0);
    signal mulr_2_28 : std_logic_vector(8 downto 0);
    signal mulr_1_29 : std_logic_vector(8 downto 0);
    signal mulr_2_29 : std_logic_vector(8 downto 0);
    signal mulr_1_30 : std_logic_vector(8 downto 0);
    signal mulr_2_30 : std_logic_vector(8 downto 0);
    signal mulr_1_31 : std_logic_vector(8 downto 0);
    signal mulr_2_31 : std_logic_vector(8 downto 0);
    signal mulr_1_32 : std_logic_vector(8 downto 0);
    signal mulr_2_32 : std_logic_vector(8 downto 0);
    signal mulr_1_33 : std_logic_vector(8 downto 0);
    signal mulr_2_33 : std_logic_vector(8 downto 0);
    signal mulr_1_34 : std_logic_vector(8 downto 0);
    signal mulr_2_34 : std_logic_vector(8 downto 0);
    signal mulr_1_35 : std_logic_vector(8 downto 0);
    signal mulr_2_35 : std_logic_vector(8 downto 0);
    signal mulr_1_36 : std_logic_vector(8 downto 0);
    signal mulr_2_36 : std_logic_vector(8 downto 0);
    signal mulr_1_37 : std_logic_vector(8 downto 0);
    signal mulr_2_37 : std_logic_vector(8 downto 0);
    signal mulr_1_38 : std_logic_vector(8 downto 0);
    signal mulr_2_38 : std_logic_vector(8 downto 0);
    signal mulr_1_39 : std_logic_vector(8 downto 0);
    signal mulr_2_39 : std_logic_vector(8 downto 0);
    signal mulr_1_40 : std_logic_vector(8 downto 0);
    signal mulr_2_40 : std_logic_vector(8 downto 0);
    signal mulr_1_41 : std_logic_vector(8 downto 0);
    signal mulr_2_41 : std_logic_vector(8 downto 0);
    signal mulr_1_42 : std_logic_vector(8 downto 0);
    signal mulr_2_42 : std_logic_vector(8 downto 0);
    signal mulr_1_43 : std_logic_vector(8 downto 0);
    signal mulr_2_43 : std_logic_vector(8 downto 0);
    signal mulr_1_44 : std_logic_vector(8 downto 0);
    signal mulr_2_44 : std_logic_vector(8 downto 0);
    signal mulr_1_45 : std_logic_vector(8 downto 0);
    signal mulr_2_45 : std_logic_vector(8 downto 0);
    signal mulr_1_46 : std_logic_vector(8 downto 0);
    signal mulr_2_46 : std_logic_vector(8 downto 0);
    signal mulr_1_47 : std_logic_vector(8 downto 0);
    signal mulr_2_47 : std_logic_vector(8 downto 0);
    signal mulr_1_48 : std_logic_vector(8 downto 0);
    signal mulr_2_48 : std_logic_vector(8 downto 0);
    signal mulr_1_49 : std_logic_vector(8 downto 0);
    signal mulr_2_49 : std_logic_vector(8 downto 0);
    signal mulr_1_50 : std_logic_vector(8 downto 0);
    signal mulr_2_50 : std_logic_vector(8 downto 0);
    signal mulr_1_51 : std_logic_vector(8 downto 0);
    signal mulr_2_51 : std_logic_vector(8 downto 0);
    signal mulr_1_52 : std_logic_vector(8 downto 0);
    signal mulr_2_52 : std_logic_vector(8 downto 0);
    signal mulr_1_53 : std_logic_vector(8 downto 0);
    signal mulr_2_53 : std_logic_vector(8 downto 0);
    signal mulr_1_54 : std_logic_vector(8 downto 0);
    signal mulr_2_54 : std_logic_vector(8 downto 0);
    signal mulr_1_55 : std_logic_vector(8 downto 0);
    signal mulr_2_55 : std_logic_vector(8 downto 0);
    signal mulr_1_56 : std_logic_vector(8 downto 0);
    signal mulr_2_56 : std_logic_vector(8 downto 0);
    signal mulr_1_57 : std_logic_vector(8 downto 0);
    signal mulr_2_57 : std_logic_vector(8 downto 0);
    signal mulr_1_58 : std_logic_vector(8 downto 0);
    signal mulr_2_58 : std_logic_vector(8 downto 0);
    signal mulr_1_59 : std_logic_vector(8 downto 0);
    signal mulr_2_59 : std_logic_vector(8 downto 0);
    signal mulr_1_60 : std_logic_vector(8 downto 0);
    signal mulr_2_60 : std_logic_vector(8 downto 0);
    signal mulr_1_61 : std_logic_vector(8 downto 0);
    signal mulr_2_61 : std_logic_vector(8 downto 0);
    signal mulr_1_62 : std_logic_vector(8 downto 0);
    signal mulr_2_62 : std_logic_vector(8 downto 0);
    signal mulr_1_63 : std_logic_vector(8 downto 0);
    signal mulr_2_63 : std_logic_vector(8 downto 0);
    signal mulr_1_64 : std_logic_vector(8 downto 0);
    signal mulr_2_64 : std_logic_vector(8 downto 0);
    signal mulr_1_65 : std_logic_vector(8 downto 0);
    signal mulr_2_65 : std_logic_vector(8 downto 0);
    signal mulr_1_66 : std_logic_vector(8 downto 0);
    signal mulr_2_66 : std_logic_vector(8 downto 0);
    signal mulr_1_67 : std_logic_vector(8 downto 0);
    signal mulr_2_67 : std_logic_vector(8 downto 0);
    signal mulr_1_68 : std_logic_vector(8 downto 0);
    signal mulr_2_68 : std_logic_vector(8 downto 0);
    signal mulr_1_69 : std_logic_vector(8 downto 0);
    signal mulr_2_69 : std_logic_vector(8 downto 0);
    signal mulr_1_70 : std_logic_vector(8 downto 0);
    signal mulr_2_70 : std_logic_vector(8 downto 0);
    signal mulr_1_71 : std_logic_vector(8 downto 0);
    signal mulr_2_71 : std_logic_vector(8 downto 0);
    signal mulr_1_72 : std_logic_vector(8 downto 0);
    signal mulr_2_72 : std_logic_vector(8 downto 0);
    signal mulr_1_73 : std_logic_vector(8 downto 0);
    signal mulr_2_73 : std_logic_vector(8 downto 0);
    signal mulr_1_74 : std_logic_vector(8 downto 0);
    signal mulr_2_74 : std_logic_vector(8 downto 0);
    signal mulr_1_75 : std_logic_vector(8 downto 0);
    signal mulr_2_75 : std_logic_vector(8 downto 0);
    signal mulr_1_76 : std_logic_vector(8 downto 0);
    signal mulr_2_76 : std_logic_vector(8 downto 0);
    signal mulr_1_77 : std_logic_vector(8 downto 0);
    signal mulr_2_77 : std_logic_vector(8 downto 0);
    signal mulr_1_78 : std_logic_vector(8 downto 0);
    signal mulr_2_78 : std_logic_vector(8 downto 0);
    signal mulr_1_79 : std_logic_vector(8 downto 0);
    signal mulr_2_79 : std_logic_vector(8 downto 0);
    signal mulr_1_80 : std_logic_vector(8 downto 0);
    signal mulr_2_80 : std_logic_vector(8 downto 0);
    signal mulr_1_81 : std_logic_vector(8 downto 0);
    signal mulr_2_81 : std_logic_vector(8 downto 0);
    signal mulr_1_82 : std_logic_vector(8 downto 0);
    signal mulr_2_82 : std_logic_vector(8 downto 0);
    signal mulr_1_83 : std_logic_vector(8 downto 0);
    signal mulr_2_83 : std_logic_vector(8 downto 0);
    signal mulr_1_84 : std_logic_vector(8 downto 0);
    signal mulr_2_84 : std_logic_vector(8 downto 0);
    signal mulr_1_85 : std_logic_vector(8 downto 0);
    signal mulr_2_85 : std_logic_vector(8 downto 0);
    signal mulr_1_86 : std_logic_vector(8 downto 0);
    signal mulr_2_86 : std_logic_vector(8 downto 0);
    signal mulr_1_87 : std_logic_vector(8 downto 0);
    signal mulr_2_87 : std_logic_vector(8 downto 0);
    signal mulr_1_88 : std_logic_vector(8 downto 0);
    signal mulr_2_88 : std_logic_vector(8 downto 0);
    signal mulr_1_89 : std_logic_vector(8 downto 0);
    signal mulr_2_89 : std_logic_vector(8 downto 0);
    signal mulr_1_90 : std_logic_vector(8 downto 0);
    signal mulr_2_90 : std_logic_vector(8 downto 0);
    signal mulr_1_91 : std_logic_vector(8 downto 0);
    signal mulr_2_91 : std_logic_vector(8 downto 0);
    signal mulr_1_92 : std_logic_vector(8 downto 0);
    signal mulr_2_92 : std_logic_vector(8 downto 0);
    signal mulr_1_93 : std_logic_vector(8 downto 0);
    signal mulr_2_93 : std_logic_vector(8 downto 0);
    signal mulr_1_94 : std_logic_vector(8 downto 0);
    signal mulr_2_94 : std_logic_vector(8 downto 0);
    signal mulr_1_95 : std_logic_vector(8 downto 0);
    signal mulr_2_95 : std_logic_vector(8 downto 0);
    signal mulr_1_96 : std_logic_vector(8 downto 0);
    signal mulr_2_96 : std_logic_vector(8 downto 0);
    signal mulr_1_97 : std_logic_vector(8 downto 0);
    signal mulr_2_97 : std_logic_vector(8 downto 0);
    signal mulr_1_98 : std_logic_vector(8 downto 0);
    signal mulr_2_98 : std_logic_vector(8 downto 0);
    signal mulr_1_99 : std_logic_vector(8 downto 0);
    signal mulr_2_99 : std_logic_vector(8 downto 0);
    signal mulr_1_100 : std_logic_vector(8 downto 0);
    signal mulr_2_100 : std_logic_vector(8 downto 0);
    signal mulr_1_101 : std_logic_vector(8 downto 0);
    signal mulr_2_101 : std_logic_vector(8 downto 0);
    signal mulr_1_102 : std_logic_vector(8 downto 0);
    signal mulr_2_102 : std_logic_vector(8 downto 0);
    signal mulr_1_103 : std_logic_vector(8 downto 0);
    signal mulr_2_103 : std_logic_vector(8 downto 0);
    signal mulr_1_104 : std_logic_vector(8 downto 0);
    signal mulr_2_104 : std_logic_vector(8 downto 0);
    signal mulr_1_105 : std_logic_vector(8 downto 0);
    signal mulr_2_105 : std_logic_vector(8 downto 0);
    signal mulr_1_106 : std_logic_vector(8 downto 0);
    signal mulr_2_106 : std_logic_vector(8 downto 0);
    signal mulr_1_107 : std_logic_vector(8 downto 0);
    signal mulr_2_107 : std_logic_vector(8 downto 0);
    signal mulr_1_108 : std_logic_vector(8 downto 0);
    signal mulr_2_108 : std_logic_vector(8 downto 0);
    signal mulr_1_109 : std_logic_vector(8 downto 0);
    signal mulr_2_109 : std_logic_vector(8 downto 0);
    signal mulr_1_110 : std_logic_vector(8 downto 0);
    signal mulr_2_110 : std_logic_vector(8 downto 0);
    signal mulr_1_111 : std_logic_vector(8 downto 0);
    signal mulr_2_111 : std_logic_vector(8 downto 0);
    signal mulr_1_112 : std_logic_vector(8 downto 0);
    signal mulr_2_112 : std_logic_vector(8 downto 0);
    signal mulr_1_113 : std_logic_vector(8 downto 0);
    signal mulr_2_113 : std_logic_vector(8 downto 0);
    signal mulr_1_114 : std_logic_vector(8 downto 0);
    signal mulr_2_114 : std_logic_vector(8 downto 0);
    signal mulr_1_115 : std_logic_vector(8 downto 0);
    signal mulr_2_115 : std_logic_vector(8 downto 0);
    signal mulr_1_116 : std_logic_vector(8 downto 0);
    signal mulr_2_116 : std_logic_vector(8 downto 0);
    signal mulr_1_117 : std_logic_vector(8 downto 0);
    signal mulr_2_117 : std_logic_vector(8 downto 0);
    signal mulr_1_118 : std_logic_vector(8 downto 0);
    signal mulr_2_118 : std_logic_vector(8 downto 0);
    signal mulr_1_119 : std_logic_vector(8 downto 0);
    signal mulr_2_119 : std_logic_vector(8 downto 0);
    signal mulr_1_120 : std_logic_vector(8 downto 0);
    signal mulr_2_120 : std_logic_vector(8 downto 0);
    signal mulr_1_121 : std_logic_vector(8 downto 0);
    signal mulr_2_121 : std_logic_vector(8 downto 0);
    signal mulr_1_122 : std_logic_vector(8 downto 0);
    signal mulr_2_122 : std_logic_vector(8 downto 0);
    signal mulr_1_123 : std_logic_vector(8 downto 0);
    signal mulr_2_123 : std_logic_vector(8 downto 0);
    signal mulr_1_124 : std_logic_vector(8 downto 0);
    signal mulr_2_124 : std_logic_vector(8 downto 0);
    signal mulr_1_125 : std_logic_vector(8 downto 0);
    signal mulr_2_125 : std_logic_vector(8 downto 0);
    signal mulr_1_126 : std_logic_vector(8 downto 0);
    signal mulr_2_126 : std_logic_vector(8 downto 0);
    signal mulr_1_127 : std_logic_vector(8 downto 0);
    signal mulr_2_127 : std_logic_vector(8 downto 0);
    signal mulr_1_128 : std_logic_vector(8 downto 0);
    signal mulr_2_128 : std_logic_vector(8 downto 0);
    signal mulr_1_129 : std_logic_vector(8 downto 0);
    signal mulr_2_129 : std_logic_vector(8 downto 0);
    signal mulr_1_130 : std_logic_vector(8 downto 0);
    signal mulr_2_130 : std_logic_vector(8 downto 0);
    signal mulr_1_131 : std_logic_vector(8 downto 0);
    signal mulr_2_131 : std_logic_vector(8 downto 0);
    signal mulr_1_132 : std_logic_vector(8 downto 0);
    signal mulr_2_132 : std_logic_vector(8 downto 0);
    signal mulr_1_133 : std_logic_vector(8 downto 0);
    signal mulr_2_133 : std_logic_vector(8 downto 0);
    signal mulr_1_134 : std_logic_vector(8 downto 0);
    signal mulr_2_134 : std_logic_vector(8 downto 0);
    signal mulr_1_135 : std_logic_vector(8 downto 0);
    signal mulr_2_135 : std_logic_vector(8 downto 0);
    signal mulr_1_136 : std_logic_vector(8 downto 0);
    signal mulr_2_136 : std_logic_vector(8 downto 0);
    signal mulr_1_137 : std_logic_vector(8 downto 0);
    signal mulr_2_137 : std_logic_vector(8 downto 0);
    signal mulr_1_138 : std_logic_vector(8 downto 0);
    signal mulr_2_138 : std_logic_vector(8 downto 0);
    signal mulr_1_139 : std_logic_vector(8 downto 0);
    signal mulr_2_139 : std_logic_vector(8 downto 0);
    signal mulr_1_140 : std_logic_vector(8 downto 0);
    signal mulr_2_140 : std_logic_vector(8 downto 0);
    signal mulr_1_141 : std_logic_vector(8 downto 0);
    signal mulr_2_141 : std_logic_vector(8 downto 0);
    signal mulr_1_142 : std_logic_vector(8 downto 0);
    signal mulr_2_142 : std_logic_vector(8 downto 0);
    signal mulr_1_143 : std_logic_vector(8 downto 0);
    signal mulr_2_143 : std_logic_vector(8 downto 0);
    signal mulr_1_144 : std_logic_vector(8 downto 0);
    signal mulr_2_144 : std_logic_vector(8 downto 0);
    signal mulr_1_145 : std_logic_vector(8 downto 0);
    signal mulr_2_145 : std_logic_vector(8 downto 0);
    signal mulr_1_146 : std_logic_vector(8 downto 0);
    signal mulr_2_146 : std_logic_vector(8 downto 0);
    signal mulr_1_147 : std_logic_vector(8 downto 0);
    signal mulr_2_147 : std_logic_vector(8 downto 0);
    signal mulr_1_148 : std_logic_vector(8 downto 0);
    signal mulr_2_148 : std_logic_vector(8 downto 0);
    signal mulr_1_149 : std_logic_vector(8 downto 0);
    signal mulr_2_149 : std_logic_vector(8 downto 0);
    signal mulr_1_150 : std_logic_vector(8 downto 0);
    signal mulr_2_150 : std_logic_vector(8 downto 0);
    signal mulr_1_151 : std_logic_vector(8 downto 0);
    signal mulr_2_151 : std_logic_vector(8 downto 0);
    signal mulr_1_152 : std_logic_vector(8 downto 0);
    signal mulr_2_152 : std_logic_vector(8 downto 0);
    signal mulr_1_153 : std_logic_vector(8 downto 0);
    signal mulr_2_153 : std_logic_vector(8 downto 0);
    signal mulr_1_154 : std_logic_vector(8 downto 0);
    signal mulr_2_154 : std_logic_vector(8 downto 0);
    signal mulr_1_155 : std_logic_vector(8 downto 0);
    signal mulr_2_155 : std_logic_vector(8 downto 0);
    signal mulr_1_156 : std_logic_vector(8 downto 0);
    signal mulr_2_156 : std_logic_vector(8 downto 0);
    signal mulr_1_157 : std_logic_vector(8 downto 0);
    signal mulr_2_157 : std_logic_vector(8 downto 0);
    signal mulr_1_158 : std_logic_vector(8 downto 0);
    signal mulr_2_158 : std_logic_vector(8 downto 0);
    signal mulr_1_159 : std_logic_vector(8 downto 0);
    signal mulr_2_159 : std_logic_vector(8 downto 0);
    signal mulr_1_160 : std_logic_vector(8 downto 0);
    signal mulr_2_160 : std_logic_vector(8 downto 0);
    signal mulr_1_161 : std_logic_vector(8 downto 0);
    signal mulr_2_161 : std_logic_vector(8 downto 0);
    signal mulr_1_162 : std_logic_vector(8 downto 0);
    signal mulr_2_162 : std_logic_vector(8 downto 0);
    signal mulr_1_163 : std_logic_vector(8 downto 0);
    signal mulr_2_163 : std_logic_vector(8 downto 0);
    signal mulr_1_164 : std_logic_vector(8 downto 0);
    signal mulr_2_164 : std_logic_vector(8 downto 0);
    signal mulr_1_165 : std_logic_vector(8 downto 0);
    signal mulr_2_165 : std_logic_vector(8 downto 0);
    signal mulr_1_166 : std_logic_vector(8 downto 0);
    signal mulr_2_166 : std_logic_vector(8 downto 0);
    signal mulr_1_167 : std_logic_vector(8 downto 0);
    signal mulr_2_167 : std_logic_vector(8 downto 0);
    signal mulr_1_168 : std_logic_vector(8 downto 0);
    signal mulr_2_168 : std_logic_vector(8 downto 0);
    signal mulr_1_169 : std_logic_vector(8 downto 0);
    signal mulr_2_169 : std_logic_vector(8 downto 0);
    signal mulr_1_170 : std_logic_vector(8 downto 0);
    signal mulr_2_170 : std_logic_vector(8 downto 0);
    signal mulr_1_171 : std_logic_vector(8 downto 0);
    signal mulr_2_171 : std_logic_vector(8 downto 0);
    signal mulr_1_172 : std_logic_vector(8 downto 0);
    signal mulr_2_172 : std_logic_vector(8 downto 0);
    signal mulr_1_173 : std_logic_vector(8 downto 0);
    signal mulr_2_173 : std_logic_vector(8 downto 0);
    signal mulr_1_174 : std_logic_vector(8 downto 0);
    signal mulr_2_174 : std_logic_vector(8 downto 0);
    signal mulr_1_175 : std_logic_vector(8 downto 0);
    signal mulr_2_175 : std_logic_vector(8 downto 0);
    signal mulr_1_176 : std_logic_vector(8 downto 0);
    signal mulr_2_176 : std_logic_vector(8 downto 0);
    signal mulr_1_177 : std_logic_vector(8 downto 0);
    signal mulr_2_177 : std_logic_vector(8 downto 0);
    signal mulr_1_178 : std_logic_vector(8 downto 0);
    signal mulr_2_178 : std_logic_vector(8 downto 0);
    signal mulr_1_179 : std_logic_vector(8 downto 0);
    signal mulr_2_179 : std_logic_vector(8 downto 0);
    signal mulr_1_180 : std_logic_vector(8 downto 0);
    signal mulr_2_180 : std_logic_vector(8 downto 0);
    signal mulr_1_181 : std_logic_vector(8 downto 0);
    signal mulr_2_181 : std_logic_vector(8 downto 0);
    signal mulr_1_182 : std_logic_vector(8 downto 0);
    signal mulr_2_182 : std_logic_vector(8 downto 0);
    signal mulr_1_183 : std_logic_vector(8 downto 0);
    signal mulr_2_183 : std_logic_vector(8 downto 0);
    signal mulr_1_184 : std_logic_vector(8 downto 0);
    signal mulr_2_184 : std_logic_vector(8 downto 0);
    signal mulr_1_185 : std_logic_vector(8 downto 0);
    signal mulr_2_185 : std_logic_vector(8 downto 0);
    signal mulr_1_186 : std_logic_vector(8 downto 0);
    signal mulr_2_186 : std_logic_vector(8 downto 0);
    signal mulr_1_187 : std_logic_vector(8 downto 0);
    signal mulr_2_187 : std_logic_vector(8 downto 0);
    signal mulr_1_188 : std_logic_vector(8 downto 0);
    signal mulr_2_188 : std_logic_vector(8 downto 0);
    signal mulr_1_189 : std_logic_vector(8 downto 0);
    signal mulr_2_189 : std_logic_vector(8 downto 0);
    signal mulr_1_190 : std_logic_vector(8 downto 0);
    signal mulr_2_190 : std_logic_vector(8 downto 0);
    signal mulr_1_191 : std_logic_vector(8 downto 0);
    signal mulr_2_191 : std_logic_vector(8 downto 0);
    signal mulr_1_192 : std_logic_vector(8 downto 0);
    signal mulr_2_192 : std_logic_vector(8 downto 0);
    signal mulr_1_193 : std_logic_vector(8 downto 0);
    signal mulr_2_193 : std_logic_vector(8 downto 0);
    signal mulr_1_194 : std_logic_vector(8 downto 0);
    signal mulr_2_194 : std_logic_vector(8 downto 0);
    signal mulr_1_195 : std_logic_vector(8 downto 0);
    signal mulr_2_195 : std_logic_vector(8 downto 0);
    signal mulr_1_196 : std_logic_vector(8 downto 0);
    signal mulr_2_196 : std_logic_vector(8 downto 0);
    signal mulr_1_197 : std_logic_vector(8 downto 0);
    signal mulr_2_197 : std_logic_vector(8 downto 0);
    signal mulr_1_198 : std_logic_vector(8 downto 0);
    signal mulr_2_198 : std_logic_vector(8 downto 0);
    signal mulr_1_199 : std_logic_vector(8 downto 0);
    signal mulr_2_199 : std_logic_vector(8 downto 0);
    signal mulr_1_200 : std_logic_vector(8 downto 0);
    signal mulr_2_200 : std_logic_vector(8 downto 0);
    signal mulr_1_201 : std_logic_vector(8 downto 0);
    signal mulr_2_201 : std_logic_vector(8 downto 0);
    signal mulr_1_202 : std_logic_vector(8 downto 0);
    signal mulr_2_202 : std_logic_vector(8 downto 0);
    signal mulr_1_203 : std_logic_vector(8 downto 0);
    signal mulr_2_203 : std_logic_vector(8 downto 0);
    signal mulr_1_204 : std_logic_vector(8 downto 0);
    signal mulr_2_204 : std_logic_vector(8 downto 0);
    signal mulr_1_205 : std_logic_vector(8 downto 0);
    signal mulr_2_205 : std_logic_vector(8 downto 0);
    signal mulr_1_206 : std_logic_vector(8 downto 0);
    signal mulr_2_206 : std_logic_vector(8 downto 0);
    signal mulr_1_207 : std_logic_vector(8 downto 0);
    signal mulr_2_207 : std_logic_vector(8 downto 0);
    signal mulr_1_208 : std_logic_vector(8 downto 0);
    signal mulr_2_208 : std_logic_vector(8 downto 0);
    signal mulr_1_209 : std_logic_vector(8 downto 0);
    signal mulr_2_209 : std_logic_vector(8 downto 0);
    signal mulr_1_210 : std_logic_vector(8 downto 0);
    signal mulr_2_210 : std_logic_vector(8 downto 0);
    signal mulr_1_211 : std_logic_vector(8 downto 0);
    signal mulr_2_211 : std_logic_vector(8 downto 0);
    signal mulr_1_212 : std_logic_vector(8 downto 0);
    signal mulr_2_212 : std_logic_vector(8 downto 0);
    signal mulr_1_213 : std_logic_vector(8 downto 0);
    signal mulr_2_213 : std_logic_vector(8 downto 0);
    signal mulr_1_214 : std_logic_vector(8 downto 0);
    signal mulr_2_214 : std_logic_vector(8 downto 0);
    signal mulr_1_215 : std_logic_vector(8 downto 0);
    signal mulr_2_215 : std_logic_vector(8 downto 0);
    signal mulr_1_216 : std_logic_vector(8 downto 0);
    signal mulr_2_216 : std_logic_vector(8 downto 0);
    signal mulr_1_217 : std_logic_vector(8 downto 0);
    signal mulr_2_217 : std_logic_vector(8 downto 0);
    signal mulr_1_218 : std_logic_vector(8 downto 0);
    signal mulr_2_218 : std_logic_vector(8 downto 0);
    signal mulr_1_219 : std_logic_vector(8 downto 0);
    signal mulr_2_219 : std_logic_vector(8 downto 0);
    signal mulr_1_220 : std_logic_vector(8 downto 0);
    signal mulr_2_220 : std_logic_vector(8 downto 0);
    signal mulr_1_221 : std_logic_vector(8 downto 0);
    signal mulr_2_221 : std_logic_vector(8 downto 0);
    signal mulr_1_222 : std_logic_vector(8 downto 0);
    signal mulr_2_222 : std_logic_vector(8 downto 0);
    signal mulr_1_223 : std_logic_vector(8 downto 0);
    signal mulr_2_223 : std_logic_vector(8 downto 0);
    signal mulr_1_224 : std_logic_vector(8 downto 0);
    signal mulr_2_224 : std_logic_vector(8 downto 0);
    signal mulr_1_225 : std_logic_vector(8 downto 0);
    signal mulr_2_225 : std_logic_vector(8 downto 0);
    signal mulr_1_226 : std_logic_vector(8 downto 0);
    signal mulr_2_226 : std_logic_vector(8 downto 0);
    signal mulr_1_227 : std_logic_vector(8 downto 0);
    signal mulr_2_227 : std_logic_vector(8 downto 0);
    signal mulr_1_228 : std_logic_vector(8 downto 0);
    signal mulr_2_228 : std_logic_vector(8 downto 0);
    signal mulr_1_229 : std_logic_vector(8 downto 0);
    signal mulr_2_229 : std_logic_vector(8 downto 0);
    signal mulr_1_230 : std_logic_vector(8 downto 0);
    signal mulr_2_230 : std_logic_vector(8 downto 0);
    signal mulr_1_231 : std_logic_vector(8 downto 0);
    signal mulr_2_231 : std_logic_vector(8 downto 0);
    signal mulr_1_232 : std_logic_vector(8 downto 0);
    signal mulr_2_232 : std_logic_vector(8 downto 0);
    signal mulr_1_233 : std_logic_vector(8 downto 0);
    signal mulr_2_233 : std_logic_vector(8 downto 0);
    signal mulr_1_234 : std_logic_vector(8 downto 0);
    signal mulr_2_234 : std_logic_vector(8 downto 0);
    signal mulr_1_235 : std_logic_vector(8 downto 0);
    signal mulr_2_235 : std_logic_vector(8 downto 0);
    signal mulr_1_236 : std_logic_vector(8 downto 0);
    signal mulr_2_236 : std_logic_vector(8 downto 0);
    signal mulr_1_237 : std_logic_vector(8 downto 0);
    signal mulr_2_237 : std_logic_vector(8 downto 0);
    signal mulr_1_238 : std_logic_vector(8 downto 0);
    signal mulr_2_238 : std_logic_vector(8 downto 0);
    signal mulr_1_239 : std_logic_vector(8 downto 0);
    signal mulr_2_239 : std_logic_vector(8 downto 0);
    signal mulr_1_240 : std_logic_vector(8 downto 0);
    signal mulr_2_240 : std_logic_vector(8 downto 0);
    signal mulr_1_241 : std_logic_vector(8 downto 0);
    signal mulr_2_241 : std_logic_vector(8 downto 0);
    signal mulr_1_242 : std_logic_vector(8 downto 0);
    signal mulr_2_242 : std_logic_vector(8 downto 0);
    signal mulr_1_243 : std_logic_vector(8 downto 0);
    signal mulr_2_243 : std_logic_vector(8 downto 0);
    signal mulr_1_244 : std_logic_vector(8 downto 0);
    signal mulr_2_244 : std_logic_vector(8 downto 0);
    signal mulr_1_245 : std_logic_vector(8 downto 0);
    signal mulr_2_245 : std_logic_vector(8 downto 0);
    signal mulr_1_246 : std_logic_vector(8 downto 0);
    signal mulr_2_246 : std_logic_vector(8 downto 0);
    signal mulr_1_247 : std_logic_vector(8 downto 0);
    signal mulr_2_247 : std_logic_vector(8 downto 0);
    signal mulr_1_248 : std_logic_vector(8 downto 0);
    signal mulr_2_248 : std_logic_vector(8 downto 0);
    signal mulr_1_249 : std_logic_vector(8 downto 0);
    signal mulr_2_249 : std_logic_vector(8 downto 0);
    signal mulr_1_250 : std_logic_vector(8 downto 0);
    signal mulr_2_250 : std_logic_vector(8 downto 0);
    signal mulr_1_251 : std_logic_vector(8 downto 0);
    signal mulr_2_251 : std_logic_vector(8 downto 0);
    signal mulr_1_252 : std_logic_vector(8 downto 0);
    signal mulr_2_252 : std_logic_vector(8 downto 0);
    signal mulr_1_253 : std_logic_vector(8 downto 0);
    signal mulr_2_253 : std_logic_vector(8 downto 0);
    signal mulr_1_254 : std_logic_vector(8 downto 0);
    signal mulr_2_254 : std_logic_vector(8 downto 0);
    signal mulr_1_255 : std_logic_vector(8 downto 0);
    signal mulr_2_255 : std_logic_vector(8 downto 0);
    signal mulr_1_256 : std_logic_vector(8 downto 0);
    signal mulr_2_256 : std_logic_vector(8 downto 0);
    signal mulr_1_257 : std_logic_vector(8 downto 0);
    signal mulr_2_257 : std_logic_vector(8 downto 0);
    signal mulr_1_258 : std_logic_vector(8 downto 0);
    signal mulr_2_258 : std_logic_vector(8 downto 0);
    signal mulr_1_259 : std_logic_vector(8 downto 0);
    signal mulr_2_259 : std_logic_vector(8 downto 0);
    signal mulr_1_260 : std_logic_vector(8 downto 0);
    signal mulr_2_260 : std_logic_vector(8 downto 0);
    signal mulr_1_261 : std_logic_vector(8 downto 0);
    signal mulr_2_261 : std_logic_vector(8 downto 0);
    signal mulr_1_262 : std_logic_vector(8 downto 0);
    signal mulr_2_262 : std_logic_vector(8 downto 0);
    signal mulr_1_263 : std_logic_vector(8 downto 0);
    signal mulr_2_263 : std_logic_vector(8 downto 0);
    signal mulr_1_264 : std_logic_vector(8 downto 0);
    signal mulr_2_264 : std_logic_vector(8 downto 0);
    signal mulr_1_265 : std_logic_vector(8 downto 0);
    signal mulr_2_265 : std_logic_vector(8 downto 0);
    signal mulr_1_266 : std_logic_vector(8 downto 0);
    signal mulr_2_266 : std_logic_vector(8 downto 0);
    signal mulr_1_267 : std_logic_vector(8 downto 0);
    signal mulr_2_267 : std_logic_vector(8 downto 0);
    signal mulr_1_268 : std_logic_vector(8 downto 0);
    signal mulr_2_268 : std_logic_vector(8 downto 0);
    signal mulr_1_269 : std_logic_vector(8 downto 0);
    signal mulr_2_269 : std_logic_vector(8 downto 0);
    signal mulr_1_270 : std_logic_vector(8 downto 0);
    signal mulr_2_270 : std_logic_vector(8 downto 0);
    signal mulr_1_271 : std_logic_vector(8 downto 0);
    signal mulr_2_271 : std_logic_vector(8 downto 0);
    signal mulr_1_272 : std_logic_vector(8 downto 0);
    signal mulr_2_272 : std_logic_vector(8 downto 0);
    signal mulr_1_273 : std_logic_vector(8 downto 0);
    signal mulr_2_273 : std_logic_vector(8 downto 0);
    signal mulr_1_274 : std_logic_vector(8 downto 0);
    signal mulr_2_274 : std_logic_vector(8 downto 0);
    signal mulr_1_275 : std_logic_vector(8 downto 0);
    signal mulr_2_275 : std_logic_vector(8 downto 0);
    signal mulr_1_276 : std_logic_vector(8 downto 0);
    signal mulr_2_276 : std_logic_vector(8 downto 0);
    signal mulr_1_277 : std_logic_vector(8 downto 0);
    signal mulr_2_277 : std_logic_vector(8 downto 0);
    signal mulr_1_278 : std_logic_vector(8 downto 0);
    signal mulr_2_278 : std_logic_vector(8 downto 0);
    signal mulr_1_279 : std_logic_vector(8 downto 0);
    signal mulr_2_279 : std_logic_vector(8 downto 0);
    signal mulr_1_280 : std_logic_vector(8 downto 0);
    signal mulr_2_280 : std_logic_vector(8 downto 0);
    signal mulr_1_281 : std_logic_vector(8 downto 0);
    signal mulr_2_281 : std_logic_vector(8 downto 0);
    signal mulr_1_282 : std_logic_vector(8 downto 0);
    signal mulr_2_282 : std_logic_vector(8 downto 0);
    signal mulr_1_283 : std_logic_vector(8 downto 0);
    signal mulr_2_283 : std_logic_vector(8 downto 0);
    signal mulr_1_284 : std_logic_vector(8 downto 0);
    signal mulr_2_284 : std_logic_vector(8 downto 0);
    signal mulr_1_285 : std_logic_vector(8 downto 0);
    signal mulr_2_285 : std_logic_vector(8 downto 0);
    signal mulr_1_286 : std_logic_vector(8 downto 0);
    signal mulr_2_286 : std_logic_vector(8 downto 0);
    signal mulr_1_287 : std_logic_vector(8 downto 0);
    signal mulr_2_287 : std_logic_vector(8 downto 0);
    signal mulr_1_288 : std_logic_vector(8 downto 0);
    signal mulr_2_288 : std_logic_vector(8 downto 0);
    signal mulr_1_289 : std_logic_vector(8 downto 0);
    signal mulr_2_289 : std_logic_vector(8 downto 0);
    signal mulr_1_290 : std_logic_vector(8 downto 0);
    signal mulr_2_290 : std_logic_vector(8 downto 0);
    signal mulr_1_291 : std_logic_vector(8 downto 0);
    signal mulr_2_291 : std_logic_vector(8 downto 0);
    signal mulr_1_292 : std_logic_vector(8 downto 0);
    signal mulr_2_292 : std_logic_vector(8 downto 0);
    signal mulr_1_293 : std_logic_vector(8 downto 0);
    signal mulr_2_293 : std_logic_vector(8 downto 0);
    signal mulr_1_294 : std_logic_vector(8 downto 0);
    signal mulr_2_294 : std_logic_vector(8 downto 0);
    signal mulr_1_295 : std_logic_vector(8 downto 0);
    signal mulr_2_295 : std_logic_vector(8 downto 0);
    signal mulr_1_296 : std_logic_vector(8 downto 0);
    signal mulr_2_296 : std_logic_vector(8 downto 0);
    signal mulr_1_297 : std_logic_vector(8 downto 0);
    signal mulr_2_297 : std_logic_vector(8 downto 0);
    signal mulr_1_298 : std_logic_vector(8 downto 0);
    signal mulr_2_298 : std_logic_vector(8 downto 0);
    signal mulr_1_299 : std_logic_vector(8 downto 0);
    signal mulr_2_299 : std_logic_vector(8 downto 0);
    signal mulr_1_300 : std_logic_vector(8 downto 0);
    signal mulr_2_300 : std_logic_vector(8 downto 0);
    signal mulr_1_301 : std_logic_vector(8 downto 0);
    signal mulr_2_301 : std_logic_vector(8 downto 0);
    signal mulr_1_302 : std_logic_vector(8 downto 0);
    signal mulr_2_302 : std_logic_vector(8 downto 0);
    signal mulr_1_303 : std_logic_vector(8 downto 0);
    signal mulr_2_303 : std_logic_vector(8 downto 0);
    signal mulr_1_304 : std_logic_vector(8 downto 0);
    signal mulr_2_304 : std_logic_vector(8 downto 0);
    signal mulr_1_305 : std_logic_vector(8 downto 0);
    signal mulr_2_305 : std_logic_vector(8 downto 0);
    signal mulr_1_306 : std_logic_vector(8 downto 0);
    signal mulr_2_306 : std_logic_vector(8 downto 0);
    signal mulr_1_307 : std_logic_vector(8 downto 0);
    signal mulr_2_307 : std_logic_vector(8 downto 0);
    signal mulr_1_308 : std_logic_vector(8 downto 0);
    signal mulr_2_308 : std_logic_vector(8 downto 0);
    signal mulr_1_309 : std_logic_vector(8 downto 0);
    signal mulr_2_309 : std_logic_vector(8 downto 0);
    signal mulr_1_310 : std_logic_vector(8 downto 0);
    signal mulr_2_310 : std_logic_vector(8 downto 0);
    signal mulr_1_311 : std_logic_vector(8 downto 0);
    signal mulr_2_311 : std_logic_vector(8 downto 0);
    signal mulr_1_312 : std_logic_vector(8 downto 0);
    signal mulr_2_312 : std_logic_vector(8 downto 0);
    signal mulr_1_313 : std_logic_vector(8 downto 0);
    signal mulr_2_313 : std_logic_vector(8 downto 0);
    signal mulr_1_314 : std_logic_vector(8 downto 0);
    signal mulr_2_314 : std_logic_vector(8 downto 0);
    signal mulr_1_315 : std_logic_vector(8 downto 0);
    signal mulr_2_315 : std_logic_vector(8 downto 0);
    signal mulr_1_316 : std_logic_vector(8 downto 0);
    signal mulr_2_316 : std_logic_vector(8 downto 0);
    signal mulr_1_317 : std_logic_vector(8 downto 0);
    signal mulr_2_317 : std_logic_vector(8 downto 0);
    signal mulr_1_318 : std_logic_vector(8 downto 0);
    signal mulr_2_318 : std_logic_vector(8 downto 0);
    signal mulr_1_319 : std_logic_vector(8 downto 0);
    signal mulr_2_319 : std_logic_vector(8 downto 0);
    signal mulr_1_320 : std_logic_vector(8 downto 0);
    signal mulr_2_320 : std_logic_vector(8 downto 0);
    signal mulr_1_321 : std_logic_vector(8 downto 0);
    signal mulr_2_321 : std_logic_vector(8 downto 0);
    signal mulr_1_322 : std_logic_vector(8 downto 0);
    signal mulr_2_322 : std_logic_vector(8 downto 0);
    signal mulr_1_323 : std_logic_vector(8 downto 0);
    signal mulr_2_323 : std_logic_vector(8 downto 0);
    signal mulr_1_324 : std_logic_vector(8 downto 0);
    signal mulr_2_324 : std_logic_vector(8 downto 0);
    signal mulr_1_325 : std_logic_vector(8 downto 0);
    signal mulr_2_325 : std_logic_vector(8 downto 0);
    signal mulr_1_326 : std_logic_vector(8 downto 0);
    signal mulr_2_326 : std_logic_vector(8 downto 0);
    signal mulr_1_327 : std_logic_vector(8 downto 0);
    signal mulr_2_327 : std_logic_vector(8 downto 0);
    signal mulr_1_328 : std_logic_vector(8 downto 0);
    signal mulr_2_328 : std_logic_vector(8 downto 0);
    signal mulr_1_329 : std_logic_vector(8 downto 0);
    signal mulr_2_329 : std_logic_vector(8 downto 0);
    signal mulr_1_330 : std_logic_vector(8 downto 0);
    signal mulr_2_330 : std_logic_vector(8 downto 0);
    signal mulr_1_331 : std_logic_vector(8 downto 0);
    signal mulr_2_331 : std_logic_vector(8 downto 0);
    signal mulr_1_332 : std_logic_vector(8 downto 0);
    signal mulr_2_332 : std_logic_vector(8 downto 0);
    signal mulr_1_333 : std_logic_vector(8 downto 0);
    signal mulr_2_333 : std_logic_vector(8 downto 0);
    signal mulr_1_334 : std_logic_vector(8 downto 0);
    signal mulr_2_334 : std_logic_vector(8 downto 0);
    signal mulr_1_335 : std_logic_vector(8 downto 0);
    signal mulr_2_335 : std_logic_vector(8 downto 0);
    signal mulr_1_336 : std_logic_vector(8 downto 0);
    signal mulr_2_336 : std_logic_vector(8 downto 0);
    signal mulr_1_337 : std_logic_vector(8 downto 0);
    signal mulr_2_337 : std_logic_vector(8 downto 0);
    signal mulr_1_338 : std_logic_vector(8 downto 0);
    signal mulr_2_338 : std_logic_vector(8 downto 0);
    signal mulr_1_339 : std_logic_vector(8 downto 0);
    signal mulr_2_339 : std_logic_vector(8 downto 0);
    signal mulr_1_340 : std_logic_vector(8 downto 0);
    signal mulr_2_340 : std_logic_vector(8 downto 0);
    signal mulr_1_341 : std_logic_vector(8 downto 0);
    signal mulr_2_341 : std_logic_vector(8 downto 0);
    signal mulr_1_342 : std_logic_vector(8 downto 0);
    signal mulr_2_342 : std_logic_vector(8 downto 0);
    signal mulr_1_343 : std_logic_vector(8 downto 0);
    signal mulr_2_343 : std_logic_vector(8 downto 0);
    signal mulr_1_344 : std_logic_vector(8 downto 0);
    signal mulr_2_344 : std_logic_vector(8 downto 0);
    signal mulr_1_345 : std_logic_vector(8 downto 0);
    signal mulr_2_345 : std_logic_vector(8 downto 0);
    signal mulr_1_346 : std_logic_vector(8 downto 0);
    signal mulr_2_346 : std_logic_vector(8 downto 0);
    signal mulr_1_347 : std_logic_vector(8 downto 0);
    signal mulr_2_347 : std_logic_vector(8 downto 0);
    signal mulr_1_348 : std_logic_vector(8 downto 0);
    signal mulr_2_348 : std_logic_vector(8 downto 0);
    signal mulr_1_349 : std_logic_vector(8 downto 0);
    signal mulr_2_349 : std_logic_vector(8 downto 0);
    signal mulr_1_350 : std_logic_vector(8 downto 0);
    signal mulr_2_350 : std_logic_vector(8 downto 0);
    signal mulr_1_351 : std_logic_vector(8 downto 0);
    signal mulr_2_351 : std_logic_vector(8 downto 0);
    signal mulr_1_352 : std_logic_vector(8 downto 0);
    signal mulr_2_352 : std_logic_vector(8 downto 0);
    signal mulr_1_353 : std_logic_vector(8 downto 0);
    signal mulr_2_353 : std_logic_vector(8 downto 0);
    signal mulr_1_354 : std_logic_vector(8 downto 0);
    signal mulr_2_354 : std_logic_vector(8 downto 0);
    signal mulr_1_355 : std_logic_vector(8 downto 0);
    signal mulr_2_355 : std_logic_vector(8 downto 0);
    signal mulr_1_356 : std_logic_vector(8 downto 0);
    signal mulr_2_356 : std_logic_vector(8 downto 0);
    signal mulr_1_357 : std_logic_vector(8 downto 0);
    signal mulr_2_357 : std_logic_vector(8 downto 0);
    signal mulr_1_358 : std_logic_vector(8 downto 0);
    signal mulr_2_358 : std_logic_vector(8 downto 0);
    signal mulr_1_359 : std_logic_vector(8 downto 0);
    signal mulr_2_359 : std_logic_vector(8 downto 0);
    signal mulr_1_360 : std_logic_vector(8 downto 0);
    signal mulr_2_360 : std_logic_vector(8 downto 0);
    signal mulr_1_361 : std_logic_vector(8 downto 0);
    signal mulr_2_361 : std_logic_vector(8 downto 0);
    signal mulr_1_362 : std_logic_vector(8 downto 0);
    signal mulr_2_362 : std_logic_vector(8 downto 0);
    signal mulr_1_363 : std_logic_vector(8 downto 0);
    signal mulr_2_363 : std_logic_vector(8 downto 0);
    signal mulr_1_364 : std_logic_vector(8 downto 0);
    signal mulr_2_364 : std_logic_vector(8 downto 0);
    signal mulr_1_365 : std_logic_vector(8 downto 0);
    signal mulr_2_365 : std_logic_vector(8 downto 0);
    signal mulr_1_366 : std_logic_vector(8 downto 0);
    signal mulr_2_366 : std_logic_vector(8 downto 0);
    signal mulr_1_367 : std_logic_vector(8 downto 0);
    signal mulr_2_367 : std_logic_vector(8 downto 0);
    signal mulr_1_368 : std_logic_vector(8 downto 0);
    signal mulr_2_368 : std_logic_vector(8 downto 0);
    signal mulr_1_369 : std_logic_vector(8 downto 0);
    signal mulr_2_369 : std_logic_vector(8 downto 0);
    signal mulr_1_370 : std_logic_vector(8 downto 0);
    signal mulr_2_370 : std_logic_vector(8 downto 0);
    signal mulr_1_371 : std_logic_vector(8 downto 0);
    signal mulr_2_371 : std_logic_vector(8 downto 0);
    signal mulr_1_372 : std_logic_vector(8 downto 0);
    signal mulr_2_372 : std_logic_vector(8 downto 0);
    signal mulr_1_373 : std_logic_vector(8 downto 0);
    signal mulr_2_373 : std_logic_vector(8 downto 0);
    signal mulr_1_374 : std_logic_vector(8 downto 0);
    signal mulr_2_374 : std_logic_vector(8 downto 0);
    signal mulr_1_375 : std_logic_vector(8 downto 0);
    signal mulr_2_375 : std_logic_vector(8 downto 0);
    signal mulr_1_376 : std_logic_vector(8 downto 0);
    signal mulr_2_376 : std_logic_vector(8 downto 0);
    signal mulr_1_377 : std_logic_vector(8 downto 0);
    signal mulr_2_377 : std_logic_vector(8 downto 0);
    signal mulr_1_378 : std_logic_vector(8 downto 0);
    signal mulr_2_378 : std_logic_vector(8 downto 0);
    signal mulr_1_379 : std_logic_vector(8 downto 0);
    signal mulr_2_379 : std_logic_vector(8 downto 0);
    signal mulr_1_380 : std_logic_vector(8 downto 0);
    signal mulr_2_380 : std_logic_vector(8 downto 0);
    signal mulr_1_381 : std_logic_vector(8 downto 0);
    signal mulr_2_381 : std_logic_vector(8 downto 0);
    signal mulr_1_382 : std_logic_vector(8 downto 0);
    signal mulr_2_382 : std_logic_vector(8 downto 0);
    signal mulr_1_383 : std_logic_vector(8 downto 0);
    signal mulr_2_383 : std_logic_vector(8 downto 0);
    signal mulr_1_384 : std_logic_vector(8 downto 0);
    signal mulr_2_384 : std_logic_vector(8 downto 0);
    signal mulr_1_385 : std_logic_vector(8 downto 0);
    signal mulr_2_385 : std_logic_vector(8 downto 0);
    signal mulr_1_386 : std_logic_vector(8 downto 0);
    signal mulr_2_386 : std_logic_vector(8 downto 0);
    signal mulr_1_387 : std_logic_vector(8 downto 0);
    signal mulr_2_387 : std_logic_vector(8 downto 0);
    signal mulr_1_388 : std_logic_vector(8 downto 0);
    signal mulr_2_388 : std_logic_vector(8 downto 0);
    signal mulr_1_389 : std_logic_vector(8 downto 0);
    signal mulr_2_389 : std_logic_vector(8 downto 0);
    signal mulr_1_390 : std_logic_vector(8 downto 0);
    signal mulr_2_390 : std_logic_vector(8 downto 0);
    signal mulr_1_391 : std_logic_vector(8 downto 0);
    signal mulr_2_391 : std_logic_vector(8 downto 0);
    signal mulr_1_392 : std_logic_vector(8 downto 0);
    signal mulr_2_392 : std_logic_vector(8 downto 0);
    signal mulr_1_393 : std_logic_vector(8 downto 0);
    signal mulr_2_393 : std_logic_vector(8 downto 0);
    signal mulr_1_394 : std_logic_vector(8 downto 0);
    signal mulr_2_394 : std_logic_vector(8 downto 0);
    signal mulr_1_395 : std_logic_vector(8 downto 0);
    signal mulr_2_395 : std_logic_vector(8 downto 0);
    signal mulr_1_396 : std_logic_vector(8 downto 0);
    signal mulr_2_396 : std_logic_vector(8 downto 0);
    signal mulr_1_397 : std_logic_vector(8 downto 0);
    signal mulr_2_397 : std_logic_vector(8 downto 0);
    signal mulr_1_398 : std_logic_vector(8 downto 0);
    signal mulr_2_398 : std_logic_vector(8 downto 0);
    signal mulr_1_399 : std_logic_vector(8 downto 0);
    signal mulr_2_399 : std_logic_vector(8 downto 0);
    signal mulr_1_400 : std_logic_vector(8 downto 0);
    signal mulr_2_400 : std_logic_vector(8 downto 0);
    signal mulr_1_401 : std_logic_vector(8 downto 0);
    signal mulr_2_401 : std_logic_vector(8 downto 0);
    signal mulr_1_402 : std_logic_vector(8 downto 0);
    signal mulr_2_402 : std_logic_vector(8 downto 0);
    signal mulr_1_403 : std_logic_vector(8 downto 0);
    signal mulr_2_403 : std_logic_vector(8 downto 0);
    signal mulr_1_404 : std_logic_vector(8 downto 0);
    signal mulr_2_404 : std_logic_vector(8 downto 0);
    signal mulr_1_405 : std_logic_vector(8 downto 0);
    signal mulr_2_405 : std_logic_vector(8 downto 0);
    signal mulr_1_406 : std_logic_vector(8 downto 0);
    signal mulr_2_406 : std_logic_vector(8 downto 0);
    signal mulr_1_407 : std_logic_vector(8 downto 0);
    signal mulr_2_407 : std_logic_vector(8 downto 0);
    signal mulr_1_408 : std_logic_vector(8 downto 0);
    signal mulr_2_408 : std_logic_vector(8 downto 0);
    signal mulr_1_409 : std_logic_vector(8 downto 0);
    signal mulr_2_409 : std_logic_vector(8 downto 0);
    signal mulr_1_410 : std_logic_vector(8 downto 0);
    signal mulr_2_410 : std_logic_vector(8 downto 0);
    signal mulr_1_411 : std_logic_vector(8 downto 0);
    signal mulr_2_411 : std_logic_vector(8 downto 0);
    signal mulr_1_412 : std_logic_vector(8 downto 0);
    signal mulr_2_412 : std_logic_vector(8 downto 0);
    signal mulr_1_413 : std_logic_vector(8 downto 0);
    signal mulr_2_413 : std_logic_vector(8 downto 0);
    signal mulr_1_414 : std_logic_vector(8 downto 0);
    signal mulr_2_414 : std_logic_vector(8 downto 0);
    signal mulr_1_415 : std_logic_vector(8 downto 0);
    signal mulr_2_415 : std_logic_vector(8 downto 0);
    signal mulr_1_416 : std_logic_vector(8 downto 0);
    signal mulr_2_416 : std_logic_vector(8 downto 0);
    signal mulr_1_417 : std_logic_vector(8 downto 0);
    signal mulr_2_417 : std_logic_vector(8 downto 0);
    signal mulr_1_418 : std_logic_vector(8 downto 0);
    signal mulr_2_418 : std_logic_vector(8 downto 0);
    signal mulr_1_419 : std_logic_vector(8 downto 0);
    signal mulr_2_419 : std_logic_vector(8 downto 0);
    signal mulr_1_420 : std_logic_vector(8 downto 0);
    signal mulr_2_420 : std_logic_vector(8 downto 0);
    signal mulr_1_421 : std_logic_vector(8 downto 0);
    signal mulr_2_421 : std_logic_vector(8 downto 0);
    signal mulr_1_422 : std_logic_vector(8 downto 0);
    signal mulr_2_422 : std_logic_vector(8 downto 0);
    signal mulr_1_423 : std_logic_vector(8 downto 0);
    signal mulr_2_423 : std_logic_vector(8 downto 0);
    signal mulr_1_424 : std_logic_vector(8 downto 0);
    signal mulr_2_424 : std_logic_vector(8 downto 0);
    signal mulr_1_425 : std_logic_vector(8 downto 0);
    signal mulr_2_425 : std_logic_vector(8 downto 0);
    signal mulr_1_426 : std_logic_vector(8 downto 0);
    signal mulr_2_426 : std_logic_vector(8 downto 0);
    signal mulr_1_427 : std_logic_vector(8 downto 0);
    signal mulr_2_427 : std_logic_vector(8 downto 0);
    signal mulr_1_428 : std_logic_vector(8 downto 0);
    signal mulr_2_428 : std_logic_vector(8 downto 0);
    signal mulr_1_429 : std_logic_vector(8 downto 0);
    signal mulr_2_429 : std_logic_vector(8 downto 0);
    signal mulr_1_430 : std_logic_vector(8 downto 0);
    signal mulr_2_430 : std_logic_vector(8 downto 0);
    signal mulr_1_431 : std_logic_vector(8 downto 0);
    signal mulr_2_431 : std_logic_vector(8 downto 0);
    signal mulr_1_432 : std_logic_vector(8 downto 0);
    signal mulr_2_432 : std_logic_vector(8 downto 0);
    signal mulr_1_433 : std_logic_vector(8 downto 0);
    signal mulr_2_433 : std_logic_vector(8 downto 0);
    signal mulr_1_434 : std_logic_vector(8 downto 0);
    signal mulr_2_434 : std_logic_vector(8 downto 0);
    signal mulr_1_435 : std_logic_vector(8 downto 0);
    signal mulr_2_435 : std_logic_vector(8 downto 0);
    signal mulr_1_436 : std_logic_vector(8 downto 0);
    signal mulr_2_436 : std_logic_vector(8 downto 0);
    signal mulr_1_437 : std_logic_vector(8 downto 0);
    signal mulr_2_437 : std_logic_vector(8 downto 0);
    signal mulr_1_438 : std_logic_vector(8 downto 0);
    signal mulr_2_438 : std_logic_vector(8 downto 0);
    signal mulr_1_439 : std_logic_vector(8 downto 0);
    signal mulr_2_439 : std_logic_vector(8 downto 0);
    signal mulr_1_440 : std_logic_vector(8 downto 0);
    signal mulr_2_440 : std_logic_vector(8 downto 0);
    signal mulr_1_441 : std_logic_vector(8 downto 0);
    signal mulr_2_441 : std_logic_vector(8 downto 0);
    signal mulr_1_442 : std_logic_vector(8 downto 0);
    signal mulr_2_442 : std_logic_vector(8 downto 0);
    signal mulr_1_443 : std_logic_vector(8 downto 0);
    signal mulr_2_443 : std_logic_vector(8 downto 0);
    signal mulr_1_444 : std_logic_vector(8 downto 0);
    signal mulr_2_444 : std_logic_vector(8 downto 0);
    signal mulr_1_445 : std_logic_vector(8 downto 0);
    signal mulr_2_445 : std_logic_vector(8 downto 0);
    signal mulr_1_446 : std_logic_vector(8 downto 0);
    signal mulr_2_446 : std_logic_vector(8 downto 0);
    signal mulr_1_447 : std_logic_vector(8 downto 0);
    signal mulr_2_447 : std_logic_vector(8 downto 0);
    signal mulr_1_448 : std_logic_vector(8 downto 0);
    signal mulr_2_448 : std_logic_vector(8 downto 0);
    signal mulr_1_449 : std_logic_vector(8 downto 0);
    signal mulr_2_449 : std_logic_vector(8 downto 0);
    signal mulr_1_450 : std_logic_vector(8 downto 0);
    signal mulr_2_450 : std_logic_vector(8 downto 0);
    signal mulr_1_451 : std_logic_vector(8 downto 0);
    signal mulr_2_451 : std_logic_vector(8 downto 0);
    signal mulr_1_452 : std_logic_vector(8 downto 0);
    signal mulr_2_452 : std_logic_vector(8 downto 0);
    signal mulr_1_453 : std_logic_vector(8 downto 0);
    signal mulr_2_453 : std_logic_vector(8 downto 0);
    signal mulr_1_454 : std_logic_vector(8 downto 0);
    signal mulr_2_454 : std_logic_vector(8 downto 0);
    signal mulr_1_455 : std_logic_vector(8 downto 0);
    signal mulr_2_455 : std_logic_vector(8 downto 0);
    signal mulr_1_456 : std_logic_vector(8 downto 0);
    signal mulr_2_456 : std_logic_vector(8 downto 0);
    signal mulr_1_457 : std_logic_vector(8 downto 0);
    signal mulr_2_457 : std_logic_vector(8 downto 0);
    signal mulr_1_458 : std_logic_vector(8 downto 0);
    signal mulr_2_458 : std_logic_vector(8 downto 0);
    signal mulr_1_459 : std_logic_vector(8 downto 0);
    signal mulr_2_459 : std_logic_vector(8 downto 0);
    signal mulr_1_460 : std_logic_vector(8 downto 0);
    signal mulr_2_460 : std_logic_vector(8 downto 0);
    signal mulr_1_461 : std_logic_vector(8 downto 0);
    signal mulr_2_461 : std_logic_vector(8 downto 0);
    signal mulr_1_462 : std_logic_vector(8 downto 0);
    signal mulr_2_462 : std_logic_vector(8 downto 0);
    signal mulr_1_463 : std_logic_vector(8 downto 0);
    signal mulr_2_463 : std_logic_vector(8 downto 0);
    signal mulr_1_464 : std_logic_vector(8 downto 0);
    signal mulr_2_464 : std_logic_vector(8 downto 0);
    signal mulr_1_465 : std_logic_vector(8 downto 0);
    signal mulr_2_465 : std_logic_vector(8 downto 0);
    signal mulr_1_466 : std_logic_vector(8 downto 0);
    signal mulr_2_466 : std_logic_vector(8 downto 0);
    signal mulr_1_467 : std_logic_vector(8 downto 0);
    signal mulr_2_467 : std_logic_vector(8 downto 0);
    signal mulr_1_468 : std_logic_vector(8 downto 0);
    signal mulr_2_468 : std_logic_vector(8 downto 0);
    signal mulr_1_469 : std_logic_vector(8 downto 0);
    signal mulr_2_469 : std_logic_vector(8 downto 0);
    signal mulr_1_470 : std_logic_vector(8 downto 0);
    signal mulr_2_470 : std_logic_vector(8 downto 0);
    signal mulr_1_471 : std_logic_vector(8 downto 0);
    signal mulr_2_471 : std_logic_vector(8 downto 0);
    signal mulr_1_472 : std_logic_vector(8 downto 0);
    signal mulr_2_472 : std_logic_vector(8 downto 0);
    signal mulr_1_473 : std_logic_vector(8 downto 0);
    signal mulr_2_473 : std_logic_vector(8 downto 0);
    signal mulr_1_474 : std_logic_vector(8 downto 0);
    signal mulr_2_474 : std_logic_vector(8 downto 0);
    signal mulr_1_475 : std_logic_vector(8 downto 0);
    signal mulr_2_475 : std_logic_vector(8 downto 0);
    signal mulr_1_476 : std_logic_vector(8 downto 0);
    signal mulr_2_476 : std_logic_vector(8 downto 0);
    signal mulr_1_477 : std_logic_vector(8 downto 0);
    signal mulr_2_477 : std_logic_vector(8 downto 0);
    signal mulr_1_478 : std_logic_vector(8 downto 0);
    signal mulr_2_478 : std_logic_vector(8 downto 0);
    signal mulr_1_479 : std_logic_vector(8 downto 0);
    signal mulr_2_479 : std_logic_vector(8 downto 0);
    signal mulr_1_480 : std_logic_vector(8 downto 0);
    signal mulr_2_480 : std_logic_vector(8 downto 0);
    signal mulr_1_481 : std_logic_vector(8 downto 0);
    signal mulr_2_481 : std_logic_vector(8 downto 0);
    signal mulr_1_482 : std_logic_vector(8 downto 0);
    signal mulr_2_482 : std_logic_vector(8 downto 0);
    signal mulr_1_483 : std_logic_vector(8 downto 0);
    signal mulr_2_483 : std_logic_vector(8 downto 0);
    signal mulr_1_484 : std_logic_vector(8 downto 0);
    signal mulr_2_484 : std_logic_vector(8 downto 0);
    signal mulr_1_485 : std_logic_vector(8 downto 0);
    signal mulr_2_485 : std_logic_vector(8 downto 0);
    signal mulr_1_486 : std_logic_vector(8 downto 0);
    signal mulr_2_486 : std_logic_vector(8 downto 0);
    signal mulr_1_487 : std_logic_vector(8 downto 0);
    signal mulr_2_487 : std_logic_vector(8 downto 0);
    signal mulr_1_488 : std_logic_vector(8 downto 0);
    signal mulr_2_488 : std_logic_vector(8 downto 0);
    signal mulr_1_489 : std_logic_vector(8 downto 0);
    signal mulr_2_489 : std_logic_vector(8 downto 0);
    signal mulr_1_490 : std_logic_vector(8 downto 0);
    signal mulr_2_490 : std_logic_vector(8 downto 0);
    signal mulr_1_491 : std_logic_vector(8 downto 0);
    signal mulr_2_491 : std_logic_vector(8 downto 0);
    signal mulr_1_492 : std_logic_vector(8 downto 0);
    signal mulr_2_492 : std_logic_vector(8 downto 0);
    signal mulr_1_493 : std_logic_vector(8 downto 0);
    signal mulr_2_493 : std_logic_vector(8 downto 0);
    signal mulr_1_494 : std_logic_vector(8 downto 0);
    signal mulr_2_494 : std_logic_vector(8 downto 0);
    signal mulr_1_495 : std_logic_vector(8 downto 0);
    signal mulr_2_495 : std_logic_vector(8 downto 0);
    signal mulr_1_496 : std_logic_vector(8 downto 0);
    signal mulr_2_496 : std_logic_vector(8 downto 0);
    signal mulr_1_497 : std_logic_vector(8 downto 0);
    signal mulr_2_497 : std_logic_vector(8 downto 0);
    signal mulr_1_498 : std_logic_vector(8 downto 0);
    signal mulr_2_498 : std_logic_vector(8 downto 0);
    signal mulr_1_499 : std_logic_vector(8 downto 0);
    signal mulr_2_499 : std_logic_vector(8 downto 0);
    signal mulr_1_500 : std_logic_vector(8 downto 0);
    signal mulr_2_500 : std_logic_vector(8 downto 0);
    signal mulr_1_501 : std_logic_vector(8 downto 0);
    signal mulr_2_501 : std_logic_vector(8 downto 0);
    signal mulr_1_502 : std_logic_vector(8 downto 0);
    signal mulr_2_502 : std_logic_vector(8 downto 0);
    signal mulr_1_503 : std_logic_vector(8 downto 0);
    signal mulr_2_503 : std_logic_vector(8 downto 0);
    signal mulr_1_504 : std_logic_vector(8 downto 0);
    signal mulr_2_504 : std_logic_vector(8 downto 0);
    signal mulr_1_505 : std_logic_vector(8 downto 0);
    signal mulr_2_505 : std_logic_vector(8 downto 0);
    signal mulr_1_506 : std_logic_vector(8 downto 0);
    signal mulr_2_506 : std_logic_vector(8 downto 0);
    signal mulr_1_507 : std_logic_vector(8 downto 0);
    signal mulr_2_507 : std_logic_vector(8 downto 0);
    signal mulr_1_508 : std_logic_vector(8 downto 0);
    signal mulr_2_508 : std_logic_vector(8 downto 0);
    signal mulr_1_509 : std_logic_vector(8 downto 0);
    signal mulr_2_509 : std_logic_vector(8 downto 0);
    signal mulr_1_510 : std_logic_vector(8 downto 0);
    signal mulr_2_510 : std_logic_vector(8 downto 0);
    signal mulr_1_511 : std_logic_vector(8 downto 0);
    signal mulr_2_511 : std_logic_vector(8 downto 0);
    signal sumr_1 : std_logic_vector(8 downto 0);
    signal sumr_2 : std_logic_vector(8 downto 0);
    signal sumr_3 : std_logic_vector(8 downto 0);
    signal sumr_4 : std_logic_vector(8 downto 0);
    signal sumr_5 : std_logic_vector(8 downto 0);
    signal sumr_6 : std_logic_vector(8 downto 0);
    signal sumr_7 : std_logic_vector(8 downto 0);
    signal sumr_8 : std_logic_vector(8 downto 0);
    signal sumr_9 : std_logic_vector(8 downto 0);
    signal sumr_10 : std_logic_vector(8 downto 0);
    signal sumr_11 : std_logic_vector(8 downto 0);
    signal sumr_12 : std_logic_vector(8 downto 0);
    signal sumr_13 : std_logic_vector(8 downto 0);
    signal sumr_14 : std_logic_vector(8 downto 0);
    signal sumr_15 : std_logic_vector(8 downto 0);
    signal sumr_16 : std_logic_vector(8 downto 0);
    signal sumr_17 : std_logic_vector(8 downto 0);
    signal sumr_18 : std_logic_vector(8 downto 0);
    signal sumr_19 : std_logic_vector(8 downto 0);
    signal sumr_20 : std_logic_vector(8 downto 0);
    signal sumr_21 : std_logic_vector(8 downto 0);
    signal sumr_22 : std_logic_vector(8 downto 0);
    signal sumr_23 : std_logic_vector(8 downto 0);
    signal sumr_24 : std_logic_vector(8 downto 0);
    signal sumr_25 : std_logic_vector(8 downto 0);
    signal sumr_26 : std_logic_vector(8 downto 0);
    signal sumr_27 : std_logic_vector(8 downto 0);
    signal sumr_28 : std_logic_vector(8 downto 0);
    signal sumr_29 : std_logic_vector(8 downto 0);
    signal sumr_30 : std_logic_vector(8 downto 0);
    signal sumr_31 : std_logic_vector(8 downto 0);
    signal sumr_32 : std_logic_vector(8 downto 0);
    signal sumr_33 : std_logic_vector(8 downto 0);
    signal sumr_34 : std_logic_vector(8 downto 0);
    signal sumr_35 : std_logic_vector(8 downto 0);
    signal sumr_36 : std_logic_vector(8 downto 0);
    signal sumr_37 : std_logic_vector(8 downto 0);
    signal sumr_38 : std_logic_vector(8 downto 0);
    signal sumr_39 : std_logic_vector(8 downto 0);
    signal sumr_40 : std_logic_vector(8 downto 0);
    signal sumr_41 : std_logic_vector(8 downto 0);
    signal sumr_42 : std_logic_vector(8 downto 0);
    signal sumr_43 : std_logic_vector(8 downto 0);
    signal sumr_44 : std_logic_vector(8 downto 0);
    signal sumr_45 : std_logic_vector(8 downto 0);
    signal sumr_46 : std_logic_vector(8 downto 0);
    signal sumr_47 : std_logic_vector(8 downto 0);
    signal sumr_48 : std_logic_vector(8 downto 0);
    signal sumr_49 : std_logic_vector(8 downto 0);
    signal sumr_50 : std_logic_vector(8 downto 0);
    signal sumr_51 : std_logic_vector(8 downto 0);
    signal sumr_52 : std_logic_vector(8 downto 0);
    signal sumr_53 : std_logic_vector(8 downto 0);
    signal sumr_54 : std_logic_vector(8 downto 0);
    signal sumr_55 : std_logic_vector(8 downto 0);
    signal sumr_56 : std_logic_vector(8 downto 0);
    signal sumr_57 : std_logic_vector(8 downto 0);
    signal sumr_58 : std_logic_vector(8 downto 0);
    signal sumr_59 : std_logic_vector(8 downto 0);
    signal sumr_60 : std_logic_vector(8 downto 0);
    signal sumr_61 : std_logic_vector(8 downto 0);
    signal sumr_62 : std_logic_vector(8 downto 0);
    signal sumr_63 : std_logic_vector(8 downto 0);
    signal sumr_64 : std_logic_vector(8 downto 0);
    signal sumr_65 : std_logic_vector(8 downto 0);
    signal sumr_66 : std_logic_vector(8 downto 0);
    signal sumr_67 : std_logic_vector(8 downto 0);
    signal sumr_68 : std_logic_vector(8 downto 0);
    signal sumr_69 : std_logic_vector(8 downto 0);
    signal sumr_70 : std_logic_vector(8 downto 0);
    signal sumr_71 : std_logic_vector(8 downto 0);
    signal sumr_72 : std_logic_vector(8 downto 0);
    signal sumr_73 : std_logic_vector(8 downto 0);
    signal sumr_74 : std_logic_vector(8 downto 0);
    signal sumr_75 : std_logic_vector(8 downto 0);
    signal sumr_76 : std_logic_vector(8 downto 0);
    signal sumr_77 : std_logic_vector(8 downto 0);
    signal sumr_78 : std_logic_vector(8 downto 0);
    signal sumr_79 : std_logic_vector(8 downto 0);
    signal sumr_80 : std_logic_vector(8 downto 0);
    signal sumr_81 : std_logic_vector(8 downto 0);
    signal sumr_82 : std_logic_vector(8 downto 0);
    signal sumr_83 : std_logic_vector(8 downto 0);
    signal sumr_84 : std_logic_vector(8 downto 0);
    signal sumr_85 : std_logic_vector(8 downto 0);
    signal sumr_86 : std_logic_vector(8 downto 0);
    signal sumr_87 : std_logic_vector(8 downto 0);
    signal sumr_88 : std_logic_vector(8 downto 0);
    signal sumr_89 : std_logic_vector(8 downto 0);
    signal sumr_90 : std_logic_vector(8 downto 0);
    signal sumr_91 : std_logic_vector(8 downto 0);
    signal sumr_92 : std_logic_vector(8 downto 0);
    signal sumr_93 : std_logic_vector(8 downto 0);
    signal sumr_94 : std_logic_vector(8 downto 0);
    signal sumr_95 : std_logic_vector(8 downto 0);
    signal sumr_96 : std_logic_vector(8 downto 0);
    signal sumr_97 : std_logic_vector(8 downto 0);
    signal sumr_98 : std_logic_vector(8 downto 0);
    signal sumr_99 : std_logic_vector(8 downto 0);
    signal sumr_100 : std_logic_vector(8 downto 0);
    signal sumr_101 : std_logic_vector(8 downto 0);
    signal sumr_102 : std_logic_vector(8 downto 0);
    signal sumr_103 : std_logic_vector(8 downto 0);
    signal sumr_104 : std_logic_vector(8 downto 0);
    signal sumr_105 : std_logic_vector(8 downto 0);
    signal sumr_106 : std_logic_vector(8 downto 0);
    signal sumr_107 : std_logic_vector(8 downto 0);
    signal sumr_108 : std_logic_vector(8 downto 0);
    signal sumr_109 : std_logic_vector(8 downto 0);
    signal sumr_110 : std_logic_vector(8 downto 0);
    signal sumr_111 : std_logic_vector(8 downto 0);
    signal sumr_112 : std_logic_vector(8 downto 0);
    signal sumr_113 : std_logic_vector(8 downto 0);
    signal sumr_114 : std_logic_vector(8 downto 0);
    signal sumr_115 : std_logic_vector(8 downto 0);
    signal sumr_116 : std_logic_vector(8 downto 0);
    signal sumr_117 : std_logic_vector(8 downto 0);
    signal sumr_118 : std_logic_vector(8 downto 0);
    signal sumr_119 : std_logic_vector(8 downto 0);
    signal sumr_120 : std_logic_vector(8 downto 0);
    signal sumr_121 : std_logic_vector(8 downto 0);
    signal sumr_122 : std_logic_vector(8 downto 0);
    signal sumr_123 : std_logic_vector(8 downto 0);
    signal sumr_124 : std_logic_vector(8 downto 0);
    signal sumr_125 : std_logic_vector(8 downto 0);
    signal sumr_126 : std_logic_vector(8 downto 0);
    signal sumr_127 : std_logic_vector(8 downto 0);
    signal sumr_128 : std_logic_vector(8 downto 0);
    signal sumr_129 : std_logic_vector(8 downto 0);
    signal sumr_130 : std_logic_vector(8 downto 0);
    signal sumr_131 : std_logic_vector(8 downto 0);
    signal sumr_132 : std_logic_vector(8 downto 0);
    signal sumr_133 : std_logic_vector(8 downto 0);
    signal sumr_134 : std_logic_vector(8 downto 0);
    signal sumr_135 : std_logic_vector(8 downto 0);
    signal sumr_136 : std_logic_vector(8 downto 0);
    signal sumr_137 : std_logic_vector(8 downto 0);
    signal sumr_138 : std_logic_vector(8 downto 0);
    signal sumr_139 : std_logic_vector(8 downto 0);
    signal sumr_140 : std_logic_vector(8 downto 0);
    signal sumr_141 : std_logic_vector(8 downto 0);
    signal sumr_142 : std_logic_vector(8 downto 0);
    signal sumr_143 : std_logic_vector(8 downto 0);
    signal sumr_144 : std_logic_vector(8 downto 0);
    signal sumr_145 : std_logic_vector(8 downto 0);
    signal sumr_146 : std_logic_vector(8 downto 0);
    signal sumr_147 : std_logic_vector(8 downto 0);
    signal sumr_148 : std_logic_vector(8 downto 0);
    signal sumr_149 : std_logic_vector(8 downto 0);
    signal sumr_150 : std_logic_vector(8 downto 0);
    signal sumr_151 : std_logic_vector(8 downto 0);
    signal sumr_152 : std_logic_vector(8 downto 0);
    signal sumr_153 : std_logic_vector(8 downto 0);
    signal sumr_154 : std_logic_vector(8 downto 0);
    signal sumr_155 : std_logic_vector(8 downto 0);
    signal sumr_156 : std_logic_vector(8 downto 0);
    signal sumr_157 : std_logic_vector(8 downto 0);
    signal sumr_158 : std_logic_vector(8 downto 0);
    signal sumr_159 : std_logic_vector(8 downto 0);
    signal sumr_160 : std_logic_vector(8 downto 0);
    signal sumr_161 : std_logic_vector(8 downto 0);
    signal sumr_162 : std_logic_vector(8 downto 0);
    signal sumr_163 : std_logic_vector(8 downto 0);
    signal sumr_164 : std_logic_vector(8 downto 0);
    signal sumr_165 : std_logic_vector(8 downto 0);
    signal sumr_166 : std_logic_vector(8 downto 0);
    signal sumr_167 : std_logic_vector(8 downto 0);
    signal sumr_168 : std_logic_vector(8 downto 0);
    signal sumr_169 : std_logic_vector(8 downto 0);
    signal sumr_170 : std_logic_vector(8 downto 0);
    signal sumr_171 : std_logic_vector(8 downto 0);
    signal sumr_172 : std_logic_vector(8 downto 0);
    signal sumr_173 : std_logic_vector(8 downto 0);
    signal sumr_174 : std_logic_vector(8 downto 0);
    signal sumr_175 : std_logic_vector(8 downto 0);
    signal sumr_176 : std_logic_vector(8 downto 0);
    signal sumr_177 : std_logic_vector(8 downto 0);
    signal sumr_178 : std_logic_vector(8 downto 0);
    signal sumr_179 : std_logic_vector(8 downto 0);
    signal sumr_180 : std_logic_vector(8 downto 0);
    signal sumr_181 : std_logic_vector(8 downto 0);
    signal sumr_182 : std_logic_vector(8 downto 0);
    signal sumr_183 : std_logic_vector(8 downto 0);
    signal sumr_184 : std_logic_vector(8 downto 0);
    signal sumr_185 : std_logic_vector(8 downto 0);
    signal sumr_186 : std_logic_vector(8 downto 0);
    signal sumr_187 : std_logic_vector(8 downto 0);
    signal sumr_188 : std_logic_vector(8 downto 0);
    signal sumr_189 : std_logic_vector(8 downto 0);
    signal sumr_190 : std_logic_vector(8 downto 0);
    signal sumr_191 : std_logic_vector(8 downto 0);
    signal sumr_192 : std_logic_vector(8 downto 0);
    signal sumr_193 : std_logic_vector(8 downto 0);
    signal sumr_194 : std_logic_vector(8 downto 0);
    signal sumr_195 : std_logic_vector(8 downto 0);
    signal sumr_196 : std_logic_vector(8 downto 0);
    signal sumr_197 : std_logic_vector(8 downto 0);
    signal sumr_198 : std_logic_vector(8 downto 0);
    signal sumr_199 : std_logic_vector(8 downto 0);
    signal sumr_200 : std_logic_vector(8 downto 0);
    signal sumr_201 : std_logic_vector(8 downto 0);
    signal sumr_202 : std_logic_vector(8 downto 0);
    signal sumr_203 : std_logic_vector(8 downto 0);
    signal sumr_204 : std_logic_vector(8 downto 0);
    signal sumr_205 : std_logic_vector(8 downto 0);
    signal sumr_206 : std_logic_vector(8 downto 0);
    signal sumr_207 : std_logic_vector(8 downto 0);
    signal sumr_208 : std_logic_vector(8 downto 0);
    signal sumr_209 : std_logic_vector(8 downto 0);
    signal sumr_210 : std_logic_vector(8 downto 0);
    signal sumr_211 : std_logic_vector(8 downto 0);
    signal sumr_212 : std_logic_vector(8 downto 0);
    signal sumr_213 : std_logic_vector(8 downto 0);
    signal sumr_214 : std_logic_vector(8 downto 0);
    signal sumr_215 : std_logic_vector(8 downto 0);
    signal sumr_216 : std_logic_vector(8 downto 0);
    signal sumr_217 : std_logic_vector(8 downto 0);
    signal sumr_218 : std_logic_vector(8 downto 0);
    signal sumr_219 : std_logic_vector(8 downto 0);
    signal sumr_220 : std_logic_vector(8 downto 0);
    signal sumr_221 : std_logic_vector(8 downto 0);
    signal sumr_222 : std_logic_vector(8 downto 0);
    signal sumr_223 : std_logic_vector(8 downto 0);
    signal sumr_224 : std_logic_vector(8 downto 0);
    signal sumr_225 : std_logic_vector(8 downto 0);
    signal sumr_226 : std_logic_vector(8 downto 0);
    signal sumr_227 : std_logic_vector(8 downto 0);
    signal sumr_228 : std_logic_vector(8 downto 0);
    signal sumr_229 : std_logic_vector(8 downto 0);
    signal sumr_230 : std_logic_vector(8 downto 0);
    signal sumr_231 : std_logic_vector(8 downto 0);
    signal sumr_232 : std_logic_vector(8 downto 0);
    signal sumr_233 : std_logic_vector(8 downto 0);
    signal sumr_234 : std_logic_vector(8 downto 0);
    signal sumr_235 : std_logic_vector(8 downto 0);
    signal sumr_236 : std_logic_vector(8 downto 0);
    signal sumr_237 : std_logic_vector(8 downto 0);
    signal sumr_238 : std_logic_vector(8 downto 0);
    signal sumr_239 : std_logic_vector(8 downto 0);
    signal sumr_240 : std_logic_vector(8 downto 0);
    signal sumr_241 : std_logic_vector(8 downto 0);
    signal sumr_242 : std_logic_vector(8 downto 0);
    signal sumr_243 : std_logic_vector(8 downto 0);
    signal sumr_244 : std_logic_vector(8 downto 0);
    signal sumr_245 : std_logic_vector(8 downto 0);
    signal sumr_246 : std_logic_vector(8 downto 0);
    signal sumr_247 : std_logic_vector(8 downto 0);
    signal sumr_248 : std_logic_vector(8 downto 0);
    signal sumr_249 : std_logic_vector(8 downto 0);
    signal sumr_250 : std_logic_vector(8 downto 0);
    signal sumr_251 : std_logic_vector(8 downto 0);
    signal sumr_252 : std_logic_vector(8 downto 0);
    signal sumr_253 : std_logic_vector(8 downto 0);
    signal sumr_254 : std_logic_vector(8 downto 0);
    signal sumr_255 : std_logic_vector(8 downto 0);
    signal sumr_256 : std_logic_vector(8 downto 0);
    signal sumr_257 : std_logic_vector(8 downto 0);
    signal sumr_258 : std_logic_vector(8 downto 0);
    signal sumr_259 : std_logic_vector(8 downto 0);
    signal sumr_260 : std_logic_vector(8 downto 0);
    signal sumr_261 : std_logic_vector(8 downto 0);
    signal sumr_262 : std_logic_vector(8 downto 0);
    signal sumr_263 : std_logic_vector(8 downto 0);
    signal sumr_264 : std_logic_vector(8 downto 0);
    signal sumr_265 : std_logic_vector(8 downto 0);
    signal sumr_266 : std_logic_vector(8 downto 0);
    signal sumr_267 : std_logic_vector(8 downto 0);
    signal sumr_268 : std_logic_vector(8 downto 0);
    signal sumr_269 : std_logic_vector(8 downto 0);
    signal sumr_270 : std_logic_vector(8 downto 0);
    signal sumr_271 : std_logic_vector(8 downto 0);
    signal sumr_272 : std_logic_vector(8 downto 0);
    signal sumr_273 : std_logic_vector(8 downto 0);
    signal sumr_274 : std_logic_vector(8 downto 0);
    signal sumr_275 : std_logic_vector(8 downto 0);
    signal sumr_276 : std_logic_vector(8 downto 0);
    signal sumr_277 : std_logic_vector(8 downto 0);
    signal sumr_278 : std_logic_vector(8 downto 0);
    signal sumr_279 : std_logic_vector(8 downto 0);
    signal sumr_280 : std_logic_vector(8 downto 0);
    signal sumr_281 : std_logic_vector(8 downto 0);
    signal sumr_282 : std_logic_vector(8 downto 0);
    signal sumr_283 : std_logic_vector(8 downto 0);
    signal sumr_284 : std_logic_vector(8 downto 0);
    signal sumr_285 : std_logic_vector(8 downto 0);
    signal sumr_286 : std_logic_vector(8 downto 0);
    signal sumr_287 : std_logic_vector(8 downto 0);
    signal sumr_288 : std_logic_vector(8 downto 0);
    signal sumr_289 : std_logic_vector(8 downto 0);
    signal sumr_290 : std_logic_vector(8 downto 0);
    signal sumr_291 : std_logic_vector(8 downto 0);
    signal sumr_292 : std_logic_vector(8 downto 0);
    signal sumr_293 : std_logic_vector(8 downto 0);
    signal sumr_294 : std_logic_vector(8 downto 0);
    signal sumr_295 : std_logic_vector(8 downto 0);
    signal sumr_296 : std_logic_vector(8 downto 0);
    signal sumr_297 : std_logic_vector(8 downto 0);
    signal sumr_298 : std_logic_vector(8 downto 0);
    signal sumr_299 : std_logic_vector(8 downto 0);
    signal sumr_300 : std_logic_vector(8 downto 0);
    signal sumr_301 : std_logic_vector(8 downto 0);
    signal sumr_302 : std_logic_vector(8 downto 0);
    signal sumr_303 : std_logic_vector(8 downto 0);
    signal sumr_304 : std_logic_vector(8 downto 0);
    signal sumr_305 : std_logic_vector(8 downto 0);
    signal sumr_306 : std_logic_vector(8 downto 0);
    signal sumr_307 : std_logic_vector(8 downto 0);
    signal sumr_308 : std_logic_vector(8 downto 0);
    signal sumr_309 : std_logic_vector(8 downto 0);
    signal sumr_310 : std_logic_vector(8 downto 0);
    signal sumr_311 : std_logic_vector(8 downto 0);
    signal sumr_312 : std_logic_vector(8 downto 0);
    signal sumr_313 : std_logic_vector(8 downto 0);
    signal sumr_314 : std_logic_vector(8 downto 0);
    signal sumr_315 : std_logic_vector(8 downto 0);
    signal sumr_316 : std_logic_vector(8 downto 0);
    signal sumr_317 : std_logic_vector(8 downto 0);
    signal sumr_318 : std_logic_vector(8 downto 0);
    signal sumr_319 : std_logic_vector(8 downto 0);
    signal sumr_320 : std_logic_vector(8 downto 0);
    signal sumr_321 : std_logic_vector(8 downto 0);
    signal sumr_322 : std_logic_vector(8 downto 0);
    signal sumr_323 : std_logic_vector(8 downto 0);
    signal sumr_324 : std_logic_vector(8 downto 0);
    signal sumr_325 : std_logic_vector(8 downto 0);
    signal sumr_326 : std_logic_vector(8 downto 0);
    signal sumr_327 : std_logic_vector(8 downto 0);
    signal sumr_328 : std_logic_vector(8 downto 0);
    signal sumr_329 : std_logic_vector(8 downto 0);
    signal sumr_330 : std_logic_vector(8 downto 0);
    signal sumr_331 : std_logic_vector(8 downto 0);
    signal sumr_332 : std_logic_vector(8 downto 0);
    signal sumr_333 : std_logic_vector(8 downto 0);
    signal sumr_334 : std_logic_vector(8 downto 0);
    signal sumr_335 : std_logic_vector(8 downto 0);
    signal sumr_336 : std_logic_vector(8 downto 0);
    signal sumr_337 : std_logic_vector(8 downto 0);
    signal sumr_338 : std_logic_vector(8 downto 0);
    signal sumr_339 : std_logic_vector(8 downto 0);
    signal sumr_340 : std_logic_vector(8 downto 0);
    signal sumr_341 : std_logic_vector(8 downto 0);
    signal sumr_342 : std_logic_vector(8 downto 0);
    signal sumr_343 : std_logic_vector(8 downto 0);
    signal sumr_344 : std_logic_vector(8 downto 0);
    signal sumr_345 : std_logic_vector(8 downto 0);
    signal sumr_346 : std_logic_vector(8 downto 0);
    signal sumr_347 : std_logic_vector(8 downto 0);
    signal sumr_348 : std_logic_vector(8 downto 0);
    signal sumr_349 : std_logic_vector(8 downto 0);
    signal sumr_350 : std_logic_vector(8 downto 0);
    signal sumr_351 : std_logic_vector(8 downto 0);
    signal sumr_352 : std_logic_vector(8 downto 0);
    signal sumr_353 : std_logic_vector(8 downto 0);
    signal sumr_354 : std_logic_vector(8 downto 0);
    signal sumr_355 : std_logic_vector(8 downto 0);
    signal sumr_356 : std_logic_vector(8 downto 0);
    signal sumr_357 : std_logic_vector(8 downto 0);
    signal sumr_358 : std_logic_vector(8 downto 0);
    signal sumr_359 : std_logic_vector(8 downto 0);
    signal sumr_360 : std_logic_vector(8 downto 0);
    signal sumr_361 : std_logic_vector(8 downto 0);
    signal sumr_362 : std_logic_vector(8 downto 0);
    signal sumr_363 : std_logic_vector(8 downto 0);
    signal sumr_364 : std_logic_vector(8 downto 0);
    signal sumr_365 : std_logic_vector(8 downto 0);
    signal sumr_366 : std_logic_vector(8 downto 0);
    signal sumr_367 : std_logic_vector(8 downto 0);
    signal sumr_368 : std_logic_vector(8 downto 0);
    signal sumr_369 : std_logic_vector(8 downto 0);
    signal sumr_370 : std_logic_vector(8 downto 0);
    signal sumr_371 : std_logic_vector(8 downto 0);
    signal sumr_372 : std_logic_vector(8 downto 0);
    signal sumr_373 : std_logic_vector(8 downto 0);
    signal sumr_374 : std_logic_vector(8 downto 0);
    signal sumr_375 : std_logic_vector(8 downto 0);
    signal sumr_376 : std_logic_vector(8 downto 0);
    signal sumr_377 : std_logic_vector(8 downto 0);
    signal sumr_378 : std_logic_vector(8 downto 0);
    signal sumr_379 : std_logic_vector(8 downto 0);
    signal sumr_380 : std_logic_vector(8 downto 0);
    signal sumr_381 : std_logic_vector(8 downto 0);
    signal sumr_382 : std_logic_vector(8 downto 0);
    signal sumr_383 : std_logic_vector(8 downto 0);
    signal sumr_384 : std_logic_vector(8 downto 0);
    signal sumr_385 : std_logic_vector(8 downto 0);
    signal sumr_386 : std_logic_vector(8 downto 0);
    signal sumr_387 : std_logic_vector(8 downto 0);
    signal sumr_388 : std_logic_vector(8 downto 0);
    signal sumr_389 : std_logic_vector(8 downto 0);
    signal sumr_390 : std_logic_vector(8 downto 0);
    signal sumr_391 : std_logic_vector(8 downto 0);
    signal sumr_392 : std_logic_vector(8 downto 0);
    signal sumr_393 : std_logic_vector(8 downto 0);
    signal sumr_394 : std_logic_vector(8 downto 0);
    signal sumr_395 : std_logic_vector(8 downto 0);
    signal sumr_396 : std_logic_vector(8 downto 0);
    signal sumr_397 : std_logic_vector(8 downto 0);
    signal sumr_398 : std_logic_vector(8 downto 0);
    signal sumr_399 : std_logic_vector(8 downto 0);
    signal sumr_400 : std_logic_vector(8 downto 0);
    signal sumr_401 : std_logic_vector(8 downto 0);
    signal sumr_402 : std_logic_vector(8 downto 0);
    signal sumr_403 : std_logic_vector(8 downto 0);
    signal sumr_404 : std_logic_vector(8 downto 0);
    signal sumr_405 : std_logic_vector(8 downto 0);
    signal sumr_406 : std_logic_vector(8 downto 0);
    signal sumr_407 : std_logic_vector(8 downto 0);
    signal sumr_408 : std_logic_vector(8 downto 0);
    signal sumr_409 : std_logic_vector(8 downto 0);
    signal sumr_410 : std_logic_vector(8 downto 0);
    signal sumr_411 : std_logic_vector(8 downto 0);
    signal sumr_412 : std_logic_vector(8 downto 0);
    signal sumr_413 : std_logic_vector(8 downto 0);
    signal sumr_414 : std_logic_vector(8 downto 0);
    signal sumr_415 : std_logic_vector(8 downto 0);
    signal sumr_416 : std_logic_vector(8 downto 0);
    signal sumr_417 : std_logic_vector(8 downto 0);
    signal sumr_418 : std_logic_vector(8 downto 0);
    signal sumr_419 : std_logic_vector(8 downto 0);
    signal sumr_420 : std_logic_vector(8 downto 0);
    signal sumr_421 : std_logic_vector(8 downto 0);
    signal sumr_422 : std_logic_vector(8 downto 0);
    signal sumr_423 : std_logic_vector(8 downto 0);
    signal sumr_424 : std_logic_vector(8 downto 0);
    signal sumr_425 : std_logic_vector(8 downto 0);
    signal sumr_426 : std_logic_vector(8 downto 0);
    signal sumr_427 : std_logic_vector(8 downto 0);
    signal sumr_428 : std_logic_vector(8 downto 0);
    signal sumr_429 : std_logic_vector(8 downto 0);
    signal sumr_430 : std_logic_vector(8 downto 0);
    signal sumr_431 : std_logic_vector(8 downto 0);
    signal sumr_432 : std_logic_vector(8 downto 0);
    signal sumr_433 : std_logic_vector(8 downto 0);
    signal sumr_434 : std_logic_vector(8 downto 0);
    signal sumr_435 : std_logic_vector(8 downto 0);
    signal sumr_436 : std_logic_vector(8 downto 0);
    signal sumr_437 : std_logic_vector(8 downto 0);
    signal sumr_438 : std_logic_vector(8 downto 0);
    signal sumr_439 : std_logic_vector(8 downto 0);
    signal sumr_440 : std_logic_vector(8 downto 0);
    signal sumr_441 : std_logic_vector(8 downto 0);
    signal sumr_442 : std_logic_vector(8 downto 0);
    signal sumr_443 : std_logic_vector(8 downto 0);
    signal sumr_444 : std_logic_vector(8 downto 0);
    signal sumr_445 : std_logic_vector(8 downto 0);
    signal sumr_446 : std_logic_vector(8 downto 0);
    signal sumr_447 : std_logic_vector(8 downto 0);
    signal sumr_448 : std_logic_vector(8 downto 0);
    signal sumr_449 : std_logic_vector(8 downto 0);
    signal sumr_450 : std_logic_vector(8 downto 0);
    signal sumr_451 : std_logic_vector(8 downto 0);
    signal sumr_452 : std_logic_vector(8 downto 0);
    signal sumr_453 : std_logic_vector(8 downto 0);
    signal sumr_454 : std_logic_vector(8 downto 0);
    signal sumr_455 : std_logic_vector(8 downto 0);
    signal sumr_456 : std_logic_vector(8 downto 0);
    signal sumr_457 : std_logic_vector(8 downto 0);
    signal sumr_458 : std_logic_vector(8 downto 0);
    signal sumr_459 : std_logic_vector(8 downto 0);
    signal sumr_460 : std_logic_vector(8 downto 0);
    signal sumr_461 : std_logic_vector(8 downto 0);
    signal sumr_462 : std_logic_vector(8 downto 0);
    signal sumr_463 : std_logic_vector(8 downto 0);
    signal sumr_464 : std_logic_vector(8 downto 0);
    signal sumr_465 : std_logic_vector(8 downto 0);
    signal sumr_466 : std_logic_vector(8 downto 0);
    signal sumr_467 : std_logic_vector(8 downto 0);
    signal sumr_468 : std_logic_vector(8 downto 0);
    signal sumr_469 : std_logic_vector(8 downto 0);
    signal sumr_470 : std_logic_vector(8 downto 0);
    signal sumr_471 : std_logic_vector(8 downto 0);
    signal sumr_472 : std_logic_vector(8 downto 0);
    signal sumr_473 : std_logic_vector(8 downto 0);
    signal sumr_474 : std_logic_vector(8 downto 0);
    signal sumr_475 : std_logic_vector(8 downto 0);
    signal sumr_476 : std_logic_vector(8 downto 0);
    signal sumr_477 : std_logic_vector(8 downto 0);
    signal sumr_478 : std_logic_vector(8 downto 0);
    signal sumr_479 : std_logic_vector(8 downto 0);
    signal sumr_480 : std_logic_vector(8 downto 0);
    signal sumr_481 : std_logic_vector(8 downto 0);
    signal sumr_482 : std_logic_vector(8 downto 0);
    signal sumr_483 : std_logic_vector(8 downto 0);
    signal sumr_484 : std_logic_vector(8 downto 0);
    signal sumr_485 : std_logic_vector(8 downto 0);
    signal sumr_486 : std_logic_vector(8 downto 0);
    signal sumr_487 : std_logic_vector(8 downto 0);
    signal sumr_488 : std_logic_vector(8 downto 0);
    signal sumr_489 : std_logic_vector(8 downto 0);
    signal sumr_490 : std_logic_vector(8 downto 0);
    signal sumr_491 : std_logic_vector(8 downto 0);
    signal sumr_492 : std_logic_vector(8 downto 0);
    signal sumr_493 : std_logic_vector(8 downto 0);
    signal sumr_494 : std_logic_vector(8 downto 0);
    signal sumr_495 : std_logic_vector(8 downto 0);
    signal sumr_496 : std_logic_vector(8 downto 0);
    signal sumr_497 : std_logic_vector(8 downto 0);
    signal sumr_498 : std_logic_vector(8 downto 0);
    signal sumr_499 : std_logic_vector(8 downto 0);
    signal sumr_500 : std_logic_vector(8 downto 0);
    signal sumr_501 : std_logic_vector(8 downto 0);
    signal sumr_502 : std_logic_vector(8 downto 0);
    signal sumr_503 : std_logic_vector(8 downto 0);
    signal sumr_504 : std_logic_vector(8 downto 0);
    signal sumr_505 : std_logic_vector(8 downto 0);
    signal sumr_506 : std_logic_vector(8 downto 0);
    signal sumr_507 : std_logic_vector(8 downto 0);
    signal sumr_508 : std_logic_vector(8 downto 0);
    signal sumr_509 : std_logic_vector(8 downto 0);
    signal sumr_510 : std_logic_vector(8 downto 0);
    signal sumr_511 : std_logic_vector(8 downto 0);
begin

mulr_1_1<=a_1;
mulc_2_1 : entity work.gfmul
port map(
a=>a_2,
b=>"000000010",
X=>mulr_2_1);

mulr_1_2<=a_1;
mulc_2_2 : entity work.gfmul
port map(
a=>a_2,
b=>"000000100",
X=>mulr_2_2);

mulr_1_3<=a_1;
mulc_2_3 : entity work.gfmul
port map(
a=>a_2,
b=>"000001000",
X=>mulr_2_3);

mulr_1_4<=a_1;
mulc_2_4 : entity work.gfmul
port map(
a=>a_2,
b=>"000010000",
X=>mulr_2_4);

mulr_1_5<=a_1;
mulc_2_5 : entity work.gfmul
port map(
a=>a_2,
b=>"000100000",
X=>mulr_2_5);

mulr_1_6<=a_1;
mulc_2_6 : entity work.gfmul
port map(
a=>a_2,
b=>"001000000",
X=>mulr_2_6);

mulr_1_7<=a_1;
mulc_2_7 : entity work.gfmul
port map(
a=>a_2,
b=>"010000000",
X=>mulr_2_7);

mulr_1_8<=a_1;
mulc_2_8 : entity work.gfmul
port map(
a=>a_2,
b=>"100000000",
X=>mulr_2_8);

mulr_1_9<=a_1;
mulc_2_9 : entity work.gfmul
port map(
a=>a_2,
b=>"000010001",
X=>mulr_2_9);

mulr_1_10<=a_1;
mulc_2_10 : entity work.gfmul
port map(
a=>a_2,
b=>"000100010",
X=>mulr_2_10);

mulr_1_11<=a_1;
mulc_2_11 : entity work.gfmul
port map(
a=>a_2,
b=>"001000100",
X=>mulr_2_11);

mulr_1_12<=a_1;
mulc_2_12 : entity work.gfmul
port map(
a=>a_2,
b=>"010001000",
X=>mulr_2_12);

mulr_1_13<=a_1;
mulc_2_13 : entity work.gfmul
port map(
a=>a_2,
b=>"100010000",
X=>mulr_2_13);

mulr_1_14<=a_1;
mulc_2_14 : entity work.gfmul
port map(
a=>a_2,
b=>"000110001",
X=>mulr_2_14);

mulr_1_15<=a_1;
mulc_2_15 : entity work.gfmul
port map(
a=>a_2,
b=>"001100010",
X=>mulr_2_15);

mulr_1_16<=a_1;
mulc_2_16 : entity work.gfmul
port map(
a=>a_2,
b=>"011000100",
X=>mulr_2_16);

mulr_1_17<=a_1;
mulc_2_17 : entity work.gfmul
port map(
a=>a_2,
b=>"110001000",
X=>mulr_2_17);

mulr_1_18<=a_1;
mulc_2_18 : entity work.gfmul
port map(
a=>a_2,
b=>"100000001",
X=>mulr_2_18);

mulr_1_19<=a_1;
mulc_2_19 : entity work.gfmul
port map(
a=>a_2,
b=>"000010011",
X=>mulr_2_19);

mulr_1_20<=a_1;
mulc_2_20 : entity work.gfmul
port map(
a=>a_2,
b=>"000100110",
X=>mulr_2_20);

mulr_1_21<=a_1;
mulc_2_21 : entity work.gfmul
port map(
a=>a_2,
b=>"001001100",
X=>mulr_2_21);

mulr_1_22<=a_1;
mulc_2_22 : entity work.gfmul
port map(
a=>a_2,
b=>"010011000",
X=>mulr_2_22);

mulr_1_23<=a_1;
mulc_2_23 : entity work.gfmul
port map(
a=>a_2,
b=>"100110000",
X=>mulr_2_23);

mulr_1_24<=a_1;
mulc_2_24 : entity work.gfmul
port map(
a=>a_2,
b=>"001110001",
X=>mulr_2_24);

mulr_1_25<=a_1;
mulc_2_25 : entity work.gfmul
port map(
a=>a_2,
b=>"011100010",
X=>mulr_2_25);

mulr_1_26<=a_1;
mulc_2_26 : entity work.gfmul
port map(
a=>a_2,
b=>"111000100",
X=>mulr_2_26);

mulr_1_27<=a_1;
mulc_2_27 : entity work.gfmul
port map(
a=>a_2,
b=>"110011001",
X=>mulr_2_27);

mulr_1_28<=a_1;
mulc_2_28 : entity work.gfmul
port map(
a=>a_2,
b=>"100100011",
X=>mulr_2_28);

mulr_1_29<=a_1;
mulc_2_29 : entity work.gfmul
port map(
a=>a_2,
b=>"001010111",
X=>mulr_2_29);

mulr_1_30<=a_1;
mulc_2_30 : entity work.gfmul
port map(
a=>a_2,
b=>"010101110",
X=>mulr_2_30);

mulr_1_31<=a_1;
mulc_2_31 : entity work.gfmul
port map(
a=>a_2,
b=>"101011100",
X=>mulr_2_31);

mulr_1_32<=a_1;
mulc_2_32 : entity work.gfmul
port map(
a=>a_2,
b=>"010101001",
X=>mulr_2_32);

mulr_1_33<=a_1;
mulc_2_33 : entity work.gfmul
port map(
a=>a_2,
b=>"101010010",
X=>mulr_2_33);

mulr_1_34<=a_1;
mulc_2_34 : entity work.gfmul
port map(
a=>a_2,
b=>"010110101",
X=>mulr_2_34);

mulr_1_35<=a_1;
mulc_2_35 : entity work.gfmul
port map(
a=>a_2,
b=>"101101010",
X=>mulr_2_35);

mulr_1_36<=a_1;
mulc_2_36 : entity work.gfmul
port map(
a=>a_2,
b=>"011000101",
X=>mulr_2_36);

mulr_1_37<=a_1;
mulc_2_37 : entity work.gfmul
port map(
a=>a_2,
b=>"110001010",
X=>mulr_2_37);

mulr_1_38<=a_1;
mulc_2_38 : entity work.gfmul
port map(
a=>a_2,
b=>"100000101",
X=>mulr_2_38);

mulr_1_39<=a_1;
mulc_2_39 : entity work.gfmul
port map(
a=>a_2,
b=>"000011011",
X=>mulr_2_39);

mulr_1_40<=a_1;
mulc_2_40 : entity work.gfmul
port map(
a=>a_2,
b=>"000110110",
X=>mulr_2_40);

mulr_1_41<=a_1;
mulc_2_41 : entity work.gfmul
port map(
a=>a_2,
b=>"001101100",
X=>mulr_2_41);

mulr_1_42<=a_1;
mulc_2_42 : entity work.gfmul
port map(
a=>a_2,
b=>"011011000",
X=>mulr_2_42);

mulr_1_43<=a_1;
mulc_2_43 : entity work.gfmul
port map(
a=>a_2,
b=>"110110000",
X=>mulr_2_43);

mulr_1_44<=a_1;
mulc_2_44 : entity work.gfmul
port map(
a=>a_2,
b=>"101110001",
X=>mulr_2_44);

mulr_1_45<=a_1;
mulc_2_45 : entity work.gfmul
port map(
a=>a_2,
b=>"011110011",
X=>mulr_2_45);

mulr_1_46<=a_1;
mulc_2_46 : entity work.gfmul
port map(
a=>a_2,
b=>"111100110",
X=>mulr_2_46);

mulr_1_47<=a_1;
mulc_2_47 : entity work.gfmul
port map(
a=>a_2,
b=>"111011101",
X=>mulr_2_47);

mulr_1_48<=a_1;
mulc_2_48 : entity work.gfmul
port map(
a=>a_2,
b=>"110101011",
X=>mulr_2_48);

mulr_1_49<=a_1;
mulc_2_49 : entity work.gfmul
port map(
a=>a_2,
b=>"101000111",
X=>mulr_2_49);

mulr_1_50<=a_1;
mulc_2_50 : entity work.gfmul
port map(
a=>a_2,
b=>"010011111",
X=>mulr_2_50);

mulr_1_51<=a_1;
mulc_2_51 : entity work.gfmul
port map(
a=>a_2,
b=>"100111110",
X=>mulr_2_51);

mulr_1_52<=a_1;
mulc_2_52 : entity work.gfmul
port map(
a=>a_2,
b=>"001101101",
X=>mulr_2_52);

mulr_1_53<=a_1;
mulc_2_53 : entity work.gfmul
port map(
a=>a_2,
b=>"011011010",
X=>mulr_2_53);

mulr_1_54<=a_1;
mulc_2_54 : entity work.gfmul
port map(
a=>a_2,
b=>"110110100",
X=>mulr_2_54);

mulr_1_55<=a_1;
mulc_2_55 : entity work.gfmul
port map(
a=>a_2,
b=>"101111001",
X=>mulr_2_55);

mulr_1_56<=a_1;
mulc_2_56 : entity work.gfmul
port map(
a=>a_2,
b=>"011100011",
X=>mulr_2_56);

mulr_1_57<=a_1;
mulc_2_57 : entity work.gfmul
port map(
a=>a_2,
b=>"111000110",
X=>mulr_2_57);

mulr_1_58<=a_1;
mulc_2_58 : entity work.gfmul
port map(
a=>a_2,
b=>"110011101",
X=>mulr_2_58);

mulr_1_59<=a_1;
mulc_2_59 : entity work.gfmul
port map(
a=>a_2,
b=>"100101011",
X=>mulr_2_59);

mulr_1_60<=a_1;
mulc_2_60 : entity work.gfmul
port map(
a=>a_2,
b=>"001000111",
X=>mulr_2_60);

mulr_1_61<=a_1;
mulc_2_61 : entity work.gfmul
port map(
a=>a_2,
b=>"010001110",
X=>mulr_2_61);

mulr_1_62<=a_1;
mulc_2_62 : entity work.gfmul
port map(
a=>a_2,
b=>"100011100",
X=>mulr_2_62);

mulr_1_63<=a_1;
mulc_2_63 : entity work.gfmul
port map(
a=>a_2,
b=>"000101001",
X=>mulr_2_63);

mulr_1_64<=a_1;
mulc_2_64 : entity work.gfmul
port map(
a=>a_2,
b=>"001010010",
X=>mulr_2_64);

mulr_1_65<=a_1;
mulc_2_65 : entity work.gfmul
port map(
a=>a_2,
b=>"010100100",
X=>mulr_2_65);

mulr_1_66<=a_1;
mulc_2_66 : entity work.gfmul
port map(
a=>a_2,
b=>"101001000",
X=>mulr_2_66);

mulr_1_67<=a_1;
mulc_2_67 : entity work.gfmul
port map(
a=>a_2,
b=>"010000001",
X=>mulr_2_67);

mulr_1_68<=a_1;
mulc_2_68 : entity work.gfmul
port map(
a=>a_2,
b=>"100000010",
X=>mulr_2_68);

mulr_1_69<=a_1;
mulc_2_69 : entity work.gfmul
port map(
a=>a_2,
b=>"000010101",
X=>mulr_2_69);

mulr_1_70<=a_1;
mulc_2_70 : entity work.gfmul
port map(
a=>a_2,
b=>"000101010",
X=>mulr_2_70);

mulr_1_71<=a_1;
mulc_2_71 : entity work.gfmul
port map(
a=>a_2,
b=>"001010100",
X=>mulr_2_71);

mulr_1_72<=a_1;
mulc_2_72 : entity work.gfmul
port map(
a=>a_2,
b=>"010101000",
X=>mulr_2_72);

mulr_1_73<=a_1;
mulc_2_73 : entity work.gfmul
port map(
a=>a_2,
b=>"101010000",
X=>mulr_2_73);

mulr_1_74<=a_1;
mulc_2_74 : entity work.gfmul
port map(
a=>a_2,
b=>"010110001",
X=>mulr_2_74);

mulr_1_75<=a_1;
mulc_2_75 : entity work.gfmul
port map(
a=>a_2,
b=>"101100010",
X=>mulr_2_75);

mulr_1_76<=a_1;
mulc_2_76 : entity work.gfmul
port map(
a=>a_2,
b=>"011010101",
X=>mulr_2_76);

mulr_1_77<=a_1;
mulc_2_77 : entity work.gfmul
port map(
a=>a_2,
b=>"110101010",
X=>mulr_2_77);

mulr_1_78<=a_1;
mulc_2_78 : entity work.gfmul
port map(
a=>a_2,
b=>"101000101",
X=>mulr_2_78);

mulr_1_79<=a_1;
mulc_2_79 : entity work.gfmul
port map(
a=>a_2,
b=>"010011011",
X=>mulr_2_79);

mulr_1_80<=a_1;
mulc_2_80 : entity work.gfmul
port map(
a=>a_2,
b=>"100110110",
X=>mulr_2_80);

mulr_1_81<=a_1;
mulc_2_81 : entity work.gfmul
port map(
a=>a_2,
b=>"001111101",
X=>mulr_2_81);

mulr_1_82<=a_1;
mulc_2_82 : entity work.gfmul
port map(
a=>a_2,
b=>"011111010",
X=>mulr_2_82);

mulr_1_83<=a_1;
mulc_2_83 : entity work.gfmul
port map(
a=>a_2,
b=>"111110100",
X=>mulr_2_83);

mulr_1_84<=a_1;
mulc_2_84 : entity work.gfmul
port map(
a=>a_2,
b=>"111111001",
X=>mulr_2_84);

mulr_1_85<=a_1;
mulc_2_85 : entity work.gfmul
port map(
a=>a_2,
b=>"111100011",
X=>mulr_2_85);

mulr_1_86<=a_1;
mulc_2_86 : entity work.gfmul
port map(
a=>a_2,
b=>"111010111",
X=>mulr_2_86);

mulr_1_87<=a_1;
mulc_2_87 : entity work.gfmul
port map(
a=>a_2,
b=>"110111111",
X=>mulr_2_87);

mulr_1_88<=a_1;
mulc_2_88 : entity work.gfmul
port map(
a=>a_2,
b=>"101101111",
X=>mulr_2_88);

mulr_1_89<=a_1;
mulc_2_89 : entity work.gfmul
port map(
a=>a_2,
b=>"011001111",
X=>mulr_2_89);

mulr_1_90<=a_1;
mulc_2_90 : entity work.gfmul
port map(
a=>a_2,
b=>"110011110",
X=>mulr_2_90);

mulr_1_91<=a_1;
mulc_2_91 : entity work.gfmul
port map(
a=>a_2,
b=>"100101101",
X=>mulr_2_91);

mulr_1_92<=a_1;
mulc_2_92 : entity work.gfmul
port map(
a=>a_2,
b=>"001001011",
X=>mulr_2_92);

mulr_1_93<=a_1;
mulc_2_93 : entity work.gfmul
port map(
a=>a_2,
b=>"010010110",
X=>mulr_2_93);

mulr_1_94<=a_1;
mulc_2_94 : entity work.gfmul
port map(
a=>a_2,
b=>"100101100",
X=>mulr_2_94);

mulr_1_95<=a_1;
mulc_2_95 : entity work.gfmul
port map(
a=>a_2,
b=>"001001001",
X=>mulr_2_95);

mulr_1_96<=a_1;
mulc_2_96 : entity work.gfmul
port map(
a=>a_2,
b=>"010010010",
X=>mulr_2_96);

mulr_1_97<=a_1;
mulc_2_97 : entity work.gfmul
port map(
a=>a_2,
b=>"100100100",
X=>mulr_2_97);

mulr_1_98<=a_1;
mulc_2_98 : entity work.gfmul
port map(
a=>a_2,
b=>"001011001",
X=>mulr_2_98);

mulr_1_99<=a_1;
mulc_2_99 : entity work.gfmul
port map(
a=>a_2,
b=>"010110010",
X=>mulr_2_99);

mulr_1_100<=a_1;
mulc_2_100 : entity work.gfmul
port map(
a=>a_2,
b=>"101100100",
X=>mulr_2_100);

mulr_1_101<=a_1;
mulc_2_101 : entity work.gfmul
port map(
a=>a_2,
b=>"011011001",
X=>mulr_2_101);

mulr_1_102<=a_1;
mulc_2_102 : entity work.gfmul
port map(
a=>a_2,
b=>"110110010",
X=>mulr_2_102);

mulr_1_103<=a_1;
mulc_2_103 : entity work.gfmul
port map(
a=>a_2,
b=>"101110101",
X=>mulr_2_103);

mulr_1_104<=a_1;
mulc_2_104 : entity work.gfmul
port map(
a=>a_2,
b=>"011111011",
X=>mulr_2_104);

mulr_1_105<=a_1;
mulc_2_105 : entity work.gfmul
port map(
a=>a_2,
b=>"111110110",
X=>mulr_2_105);

mulr_1_106<=a_1;
mulc_2_106 : entity work.gfmul
port map(
a=>a_2,
b=>"111111101",
X=>mulr_2_106);

mulr_1_107<=a_1;
mulc_2_107 : entity work.gfmul
port map(
a=>a_2,
b=>"111101011",
X=>mulr_2_107);

mulr_1_108<=a_1;
mulc_2_108 : entity work.gfmul
port map(
a=>a_2,
b=>"111000111",
X=>mulr_2_108);

mulr_1_109<=a_1;
mulc_2_109 : entity work.gfmul
port map(
a=>a_2,
b=>"110011111",
X=>mulr_2_109);

mulr_1_110<=a_1;
mulc_2_110 : entity work.gfmul
port map(
a=>a_2,
b=>"100101111",
X=>mulr_2_110);

mulr_1_111<=a_1;
mulc_2_111 : entity work.gfmul
port map(
a=>a_2,
b=>"001001111",
X=>mulr_2_111);

mulr_1_112<=a_1;
mulc_2_112 : entity work.gfmul
port map(
a=>a_2,
b=>"010011110",
X=>mulr_2_112);

mulr_1_113<=a_1;
mulc_2_113 : entity work.gfmul
port map(
a=>a_2,
b=>"100111100",
X=>mulr_2_113);

mulr_1_114<=a_1;
mulc_2_114 : entity work.gfmul
port map(
a=>a_2,
b=>"001101001",
X=>mulr_2_114);

mulr_1_115<=a_1;
mulc_2_115 : entity work.gfmul
port map(
a=>a_2,
b=>"011010010",
X=>mulr_2_115);

mulr_1_116<=a_1;
mulc_2_116 : entity work.gfmul
port map(
a=>a_2,
b=>"110100100",
X=>mulr_2_116);

mulr_1_117<=a_1;
mulc_2_117 : entity work.gfmul
port map(
a=>a_2,
b=>"101011001",
X=>mulr_2_117);

mulr_1_118<=a_1;
mulc_2_118 : entity work.gfmul
port map(
a=>a_2,
b=>"010100011",
X=>mulr_2_118);

mulr_1_119<=a_1;
mulc_2_119 : entity work.gfmul
port map(
a=>a_2,
b=>"101000110",
X=>mulr_2_119);

mulr_1_120<=a_1;
mulc_2_120 : entity work.gfmul
port map(
a=>a_2,
b=>"010011101",
X=>mulr_2_120);

mulr_1_121<=a_1;
mulc_2_121 : entity work.gfmul
port map(
a=>a_2,
b=>"100111010",
X=>mulr_2_121);

mulr_1_122<=a_1;
mulc_2_122 : entity work.gfmul
port map(
a=>a_2,
b=>"001100101",
X=>mulr_2_122);

mulr_1_123<=a_1;
mulc_2_123 : entity work.gfmul
port map(
a=>a_2,
b=>"011001010",
X=>mulr_2_123);

mulr_1_124<=a_1;
mulc_2_124 : entity work.gfmul
port map(
a=>a_2,
b=>"110010100",
X=>mulr_2_124);

mulr_1_125<=a_1;
mulc_2_125 : entity work.gfmul
port map(
a=>a_2,
b=>"100111001",
X=>mulr_2_125);

mulr_1_126<=a_1;
mulc_2_126 : entity work.gfmul
port map(
a=>a_2,
b=>"001100011",
X=>mulr_2_126);

mulr_1_127<=a_1;
mulc_2_127 : entity work.gfmul
port map(
a=>a_2,
b=>"011000110",
X=>mulr_2_127);

mulr_1_128<=a_1;
mulc_2_128 : entity work.gfmul
port map(
a=>a_2,
b=>"110001100",
X=>mulr_2_128);

mulr_1_129<=a_1;
mulc_2_129 : entity work.gfmul
port map(
a=>a_2,
b=>"100001001",
X=>mulr_2_129);

mulr_1_130<=a_1;
mulc_2_130 : entity work.gfmul
port map(
a=>a_2,
b=>"000000011",
X=>mulr_2_130);

mulr_1_131<=a_1;
mulc_2_131 : entity work.gfmul
port map(
a=>a_2,
b=>"000000110",
X=>mulr_2_131);

mulr_1_132<=a_1;
mulc_2_132 : entity work.gfmul
port map(
a=>a_2,
b=>"000001100",
X=>mulr_2_132);

mulr_1_133<=a_1;
mulc_2_133 : entity work.gfmul
port map(
a=>a_2,
b=>"000011000",
X=>mulr_2_133);

mulr_1_134<=a_1;
mulc_2_134 : entity work.gfmul
port map(
a=>a_2,
b=>"000110000",
X=>mulr_2_134);

mulr_1_135<=a_1;
mulc_2_135 : entity work.gfmul
port map(
a=>a_2,
b=>"001100000",
X=>mulr_2_135);

mulr_1_136<=a_1;
mulc_2_136 : entity work.gfmul
port map(
a=>a_2,
b=>"011000000",
X=>mulr_2_136);

mulr_1_137<=a_1;
mulc_2_137 : entity work.gfmul
port map(
a=>a_2,
b=>"110000000",
X=>mulr_2_137);

mulr_1_138<=a_1;
mulc_2_138 : entity work.gfmul
port map(
a=>a_2,
b=>"100010001",
X=>mulr_2_138);

mulr_1_139<=a_1;
mulc_2_139 : entity work.gfmul
port map(
a=>a_2,
b=>"000110011",
X=>mulr_2_139);

mulr_1_140<=a_1;
mulc_2_140 : entity work.gfmul
port map(
a=>a_2,
b=>"001100110",
X=>mulr_2_140);

mulr_1_141<=a_1;
mulc_2_141 : entity work.gfmul
port map(
a=>a_2,
b=>"011001100",
X=>mulr_2_141);

mulr_1_142<=a_1;
mulc_2_142 : entity work.gfmul
port map(
a=>a_2,
b=>"110011000",
X=>mulr_2_142);

mulr_1_143<=a_1;
mulc_2_143 : entity work.gfmul
port map(
a=>a_2,
b=>"100100001",
X=>mulr_2_143);

mulr_1_144<=a_1;
mulc_2_144 : entity work.gfmul
port map(
a=>a_2,
b=>"001010011",
X=>mulr_2_144);

mulr_1_145<=a_1;
mulc_2_145 : entity work.gfmul
port map(
a=>a_2,
b=>"010100110",
X=>mulr_2_145);

mulr_1_146<=a_1;
mulc_2_146 : entity work.gfmul
port map(
a=>a_2,
b=>"101001100",
X=>mulr_2_146);

mulr_1_147<=a_1;
mulc_2_147 : entity work.gfmul
port map(
a=>a_2,
b=>"010001001",
X=>mulr_2_147);

mulr_1_148<=a_1;
mulc_2_148 : entity work.gfmul
port map(
a=>a_2,
b=>"100010010",
X=>mulr_2_148);

mulr_1_149<=a_1;
mulc_2_149 : entity work.gfmul
port map(
a=>a_2,
b=>"000110101",
X=>mulr_2_149);

mulr_1_150<=a_1;
mulc_2_150 : entity work.gfmul
port map(
a=>a_2,
b=>"001101010",
X=>mulr_2_150);

mulr_1_151<=a_1;
mulc_2_151 : entity work.gfmul
port map(
a=>a_2,
b=>"011010100",
X=>mulr_2_151);

mulr_1_152<=a_1;
mulc_2_152 : entity work.gfmul
port map(
a=>a_2,
b=>"110101000",
X=>mulr_2_152);

mulr_1_153<=a_1;
mulc_2_153 : entity work.gfmul
port map(
a=>a_2,
b=>"101000001",
X=>mulr_2_153);

mulr_1_154<=a_1;
mulc_2_154 : entity work.gfmul
port map(
a=>a_2,
b=>"010010011",
X=>mulr_2_154);

mulr_1_155<=a_1;
mulc_2_155 : entity work.gfmul
port map(
a=>a_2,
b=>"100100110",
X=>mulr_2_155);

mulr_1_156<=a_1;
mulc_2_156 : entity work.gfmul
port map(
a=>a_2,
b=>"001011101",
X=>mulr_2_156);

mulr_1_157<=a_1;
mulc_2_157 : entity work.gfmul
port map(
a=>a_2,
b=>"010111010",
X=>mulr_2_157);

mulr_1_158<=a_1;
mulc_2_158 : entity work.gfmul
port map(
a=>a_2,
b=>"101110100",
X=>mulr_2_158);

mulr_1_159<=a_1;
mulc_2_159 : entity work.gfmul
port map(
a=>a_2,
b=>"011111001",
X=>mulr_2_159);

mulr_1_160<=a_1;
mulc_2_160 : entity work.gfmul
port map(
a=>a_2,
b=>"111110010",
X=>mulr_2_160);

mulr_1_161<=a_1;
mulc_2_161 : entity work.gfmul
port map(
a=>a_2,
b=>"111110101",
X=>mulr_2_161);

mulr_1_162<=a_1;
mulc_2_162 : entity work.gfmul
port map(
a=>a_2,
b=>"111111011",
X=>mulr_2_162);

mulr_1_163<=a_1;
mulc_2_163 : entity work.gfmul
port map(
a=>a_2,
b=>"111100111",
X=>mulr_2_163);

mulr_1_164<=a_1;
mulc_2_164 : entity work.gfmul
port map(
a=>a_2,
b=>"111011111",
X=>mulr_2_164);

mulr_1_165<=a_1;
mulc_2_165 : entity work.gfmul
port map(
a=>a_2,
b=>"110101111",
X=>mulr_2_165);

mulr_1_166<=a_1;
mulc_2_166 : entity work.gfmul
port map(
a=>a_2,
b=>"101001111",
X=>mulr_2_166);

mulr_1_167<=a_1;
mulc_2_167 : entity work.gfmul
port map(
a=>a_2,
b=>"010001111",
X=>mulr_2_167);

mulr_1_168<=a_1;
mulc_2_168 : entity work.gfmul
port map(
a=>a_2,
b=>"100011110",
X=>mulr_2_168);

mulr_1_169<=a_1;
mulc_2_169 : entity work.gfmul
port map(
a=>a_2,
b=>"000101101",
X=>mulr_2_169);

mulr_1_170<=a_1;
mulc_2_170 : entity work.gfmul
port map(
a=>a_2,
b=>"001011010",
X=>mulr_2_170);

mulr_1_171<=a_1;
mulc_2_171 : entity work.gfmul
port map(
a=>a_2,
b=>"010110100",
X=>mulr_2_171);

mulr_1_172<=a_1;
mulc_2_172 : entity work.gfmul
port map(
a=>a_2,
b=>"101101000",
X=>mulr_2_172);

mulr_1_173<=a_1;
mulc_2_173 : entity work.gfmul
port map(
a=>a_2,
b=>"011000001",
X=>mulr_2_173);

mulr_1_174<=a_1;
mulc_2_174 : entity work.gfmul
port map(
a=>a_2,
b=>"110000010",
X=>mulr_2_174);

mulr_1_175<=a_1;
mulc_2_175 : entity work.gfmul
port map(
a=>a_2,
b=>"100010101",
X=>mulr_2_175);

mulr_1_176<=a_1;
mulc_2_176 : entity work.gfmul
port map(
a=>a_2,
b=>"000111011",
X=>mulr_2_176);

mulr_1_177<=a_1;
mulc_2_177 : entity work.gfmul
port map(
a=>a_2,
b=>"001110110",
X=>mulr_2_177);

mulr_1_178<=a_1;
mulc_2_178 : entity work.gfmul
port map(
a=>a_2,
b=>"011101100",
X=>mulr_2_178);

mulr_1_179<=a_1;
mulc_2_179 : entity work.gfmul
port map(
a=>a_2,
b=>"111011000",
X=>mulr_2_179);

mulr_1_180<=a_1;
mulc_2_180 : entity work.gfmul
port map(
a=>a_2,
b=>"110100001",
X=>mulr_2_180);

mulr_1_181<=a_1;
mulc_2_181 : entity work.gfmul
port map(
a=>a_2,
b=>"101010011",
X=>mulr_2_181);

mulr_1_182<=a_1;
mulc_2_182 : entity work.gfmul
port map(
a=>a_2,
b=>"010110111",
X=>mulr_2_182);

mulr_1_183<=a_1;
mulc_2_183 : entity work.gfmul
port map(
a=>a_2,
b=>"101101110",
X=>mulr_2_183);

mulr_1_184<=a_1;
mulc_2_184 : entity work.gfmul
port map(
a=>a_2,
b=>"011001101",
X=>mulr_2_184);

mulr_1_185<=a_1;
mulc_2_185 : entity work.gfmul
port map(
a=>a_2,
b=>"110011010",
X=>mulr_2_185);

mulr_1_186<=a_1;
mulc_2_186 : entity work.gfmul
port map(
a=>a_2,
b=>"100100101",
X=>mulr_2_186);

mulr_1_187<=a_1;
mulc_2_187 : entity work.gfmul
port map(
a=>a_2,
b=>"001011011",
X=>mulr_2_187);

mulr_1_188<=a_1;
mulc_2_188 : entity work.gfmul
port map(
a=>a_2,
b=>"010110110",
X=>mulr_2_188);

mulr_1_189<=a_1;
mulc_2_189 : entity work.gfmul
port map(
a=>a_2,
b=>"101101100",
X=>mulr_2_189);

mulr_1_190<=a_1;
mulc_2_190 : entity work.gfmul
port map(
a=>a_2,
b=>"011001001",
X=>mulr_2_190);

mulr_1_191<=a_1;
mulc_2_191 : entity work.gfmul
port map(
a=>a_2,
b=>"110010010",
X=>mulr_2_191);

mulr_1_192<=a_1;
mulc_2_192 : entity work.gfmul
port map(
a=>a_2,
b=>"100110101",
X=>mulr_2_192);

mulr_1_193<=a_1;
mulc_2_193 : entity work.gfmul
port map(
a=>a_2,
b=>"001111011",
X=>mulr_2_193);

mulr_1_194<=a_1;
mulc_2_194 : entity work.gfmul
port map(
a=>a_2,
b=>"011110110",
X=>mulr_2_194);

mulr_1_195<=a_1;
mulc_2_195 : entity work.gfmul
port map(
a=>a_2,
b=>"111101100",
X=>mulr_2_195);

mulr_1_196<=a_1;
mulc_2_196 : entity work.gfmul
port map(
a=>a_2,
b=>"111001001",
X=>mulr_2_196);

mulr_1_197<=a_1;
mulc_2_197 : entity work.gfmul
port map(
a=>a_2,
b=>"110000011",
X=>mulr_2_197);

mulr_1_198<=a_1;
mulc_2_198 : entity work.gfmul
port map(
a=>a_2,
b=>"100010111",
X=>mulr_2_198);

mulr_1_199<=a_1;
mulc_2_199 : entity work.gfmul
port map(
a=>a_2,
b=>"000111111",
X=>mulr_2_199);

mulr_1_200<=a_1;
mulc_2_200 : entity work.gfmul
port map(
a=>a_2,
b=>"001111110",
X=>mulr_2_200);

mulr_1_201<=a_1;
mulc_2_201 : entity work.gfmul
port map(
a=>a_2,
b=>"011111100",
X=>mulr_2_201);

mulr_1_202<=a_1;
mulc_2_202 : entity work.gfmul
port map(
a=>a_2,
b=>"111111000",
X=>mulr_2_202);

mulr_1_203<=a_1;
mulc_2_203 : entity work.gfmul
port map(
a=>a_2,
b=>"111100001",
X=>mulr_2_203);

mulr_1_204<=a_1;
mulc_2_204 : entity work.gfmul
port map(
a=>a_2,
b=>"111010011",
X=>mulr_2_204);

mulr_1_205<=a_1;
mulc_2_205 : entity work.gfmul
port map(
a=>a_2,
b=>"110110111",
X=>mulr_2_205);

mulr_1_206<=a_1;
mulc_2_206 : entity work.gfmul
port map(
a=>a_2,
b=>"101111111",
X=>mulr_2_206);

mulr_1_207<=a_1;
mulc_2_207 : entity work.gfmul
port map(
a=>a_2,
b=>"011101111",
X=>mulr_2_207);

mulr_1_208<=a_1;
mulc_2_208 : entity work.gfmul
port map(
a=>a_2,
b=>"111011110",
X=>mulr_2_208);

mulr_1_209<=a_1;
mulc_2_209 : entity work.gfmul
port map(
a=>a_2,
b=>"110101101",
X=>mulr_2_209);

mulr_1_210<=a_1;
mulc_2_210 : entity work.gfmul
port map(
a=>a_2,
b=>"101001011",
X=>mulr_2_210);

mulr_1_211<=a_1;
mulc_2_211 : entity work.gfmul
port map(
a=>a_2,
b=>"010000111",
X=>mulr_2_211);

mulr_1_212<=a_1;
mulc_2_212 : entity work.gfmul
port map(
a=>a_2,
b=>"100001110",
X=>mulr_2_212);

mulr_1_213<=a_1;
mulc_2_213 : entity work.gfmul
port map(
a=>a_2,
b=>"000001101",
X=>mulr_2_213);

mulr_1_214<=a_1;
mulc_2_214 : entity work.gfmul
port map(
a=>a_2,
b=>"000011010",
X=>mulr_2_214);

mulr_1_215<=a_1;
mulc_2_215 : entity work.gfmul
port map(
a=>a_2,
b=>"000110100",
X=>mulr_2_215);

mulr_1_216<=a_1;
mulc_2_216 : entity work.gfmul
port map(
a=>a_2,
b=>"001101000",
X=>mulr_2_216);

mulr_1_217<=a_1;
mulc_2_217 : entity work.gfmul
port map(
a=>a_2,
b=>"011010000",
X=>mulr_2_217);

mulr_1_218<=a_1;
mulc_2_218 : entity work.gfmul
port map(
a=>a_2,
b=>"110100000",
X=>mulr_2_218);

mulr_1_219<=a_1;
mulc_2_219 : entity work.gfmul
port map(
a=>a_2,
b=>"101010001",
X=>mulr_2_219);

mulr_1_220<=a_1;
mulc_2_220 : entity work.gfmul
port map(
a=>a_2,
b=>"010110011",
X=>mulr_2_220);

mulr_1_221<=a_1;
mulc_2_221 : entity work.gfmul
port map(
a=>a_2,
b=>"101100110",
X=>mulr_2_221);

mulr_1_222<=a_1;
mulc_2_222 : entity work.gfmul
port map(
a=>a_2,
b=>"011011101",
X=>mulr_2_222);

mulr_1_223<=a_1;
mulc_2_223 : entity work.gfmul
port map(
a=>a_2,
b=>"110111010",
X=>mulr_2_223);

mulr_1_224<=a_1;
mulc_2_224 : entity work.gfmul
port map(
a=>a_2,
b=>"101100101",
X=>mulr_2_224);

mulr_1_225<=a_1;
mulc_2_225 : entity work.gfmul
port map(
a=>a_2,
b=>"011011011",
X=>mulr_2_225);

mulr_1_226<=a_1;
mulc_2_226 : entity work.gfmul
port map(
a=>a_2,
b=>"110110110",
X=>mulr_2_226);

mulr_1_227<=a_1;
mulc_2_227 : entity work.gfmul
port map(
a=>a_2,
b=>"101111101",
X=>mulr_2_227);

mulr_1_228<=a_1;
mulc_2_228 : entity work.gfmul
port map(
a=>a_2,
b=>"011101011",
X=>mulr_2_228);

mulr_1_229<=a_1;
mulc_2_229 : entity work.gfmul
port map(
a=>a_2,
b=>"111010110",
X=>mulr_2_229);

mulr_1_230<=a_1;
mulc_2_230 : entity work.gfmul
port map(
a=>a_2,
b=>"110111101",
X=>mulr_2_230);

mulr_1_231<=a_1;
mulc_2_231 : entity work.gfmul
port map(
a=>a_2,
b=>"101101011",
X=>mulr_2_231);

mulr_1_232<=a_1;
mulc_2_232 : entity work.gfmul
port map(
a=>a_2,
b=>"011000111",
X=>mulr_2_232);

mulr_1_233<=a_1;
mulc_2_233 : entity work.gfmul
port map(
a=>a_2,
b=>"110001110",
X=>mulr_2_233);

mulr_1_234<=a_1;
mulc_2_234 : entity work.gfmul
port map(
a=>a_2,
b=>"100001101",
X=>mulr_2_234);

mulr_1_235<=a_1;
mulc_2_235 : entity work.gfmul
port map(
a=>a_2,
b=>"000001011",
X=>mulr_2_235);

mulr_1_236<=a_1;
mulc_2_236 : entity work.gfmul
port map(
a=>a_2,
b=>"000010110",
X=>mulr_2_236);

mulr_1_237<=a_1;
mulc_2_237 : entity work.gfmul
port map(
a=>a_2,
b=>"000101100",
X=>mulr_2_237);

mulr_1_238<=a_1;
mulc_2_238 : entity work.gfmul
port map(
a=>a_2,
b=>"001011000",
X=>mulr_2_238);

mulr_1_239<=a_1;
mulc_2_239 : entity work.gfmul
port map(
a=>a_2,
b=>"010110000",
X=>mulr_2_239);

mulr_1_240<=a_1;
mulc_2_240 : entity work.gfmul
port map(
a=>a_2,
b=>"101100000",
X=>mulr_2_240);

mulr_1_241<=a_1;
mulc_2_241 : entity work.gfmul
port map(
a=>a_2,
b=>"011010001",
X=>mulr_2_241);

mulr_1_242<=a_1;
mulc_2_242 : entity work.gfmul
port map(
a=>a_2,
b=>"110100010",
X=>mulr_2_242);

mulr_1_243<=a_1;
mulc_2_243 : entity work.gfmul
port map(
a=>a_2,
b=>"101010101",
X=>mulr_2_243);

mulr_1_244<=a_1;
mulc_2_244 : entity work.gfmul
port map(
a=>a_2,
b=>"010111011",
X=>mulr_2_244);

mulr_1_245<=a_1;
mulc_2_245 : entity work.gfmul
port map(
a=>a_2,
b=>"101110110",
X=>mulr_2_245);

mulr_1_246<=a_1;
mulc_2_246 : entity work.gfmul
port map(
a=>a_2,
b=>"011111101",
X=>mulr_2_246);

mulr_1_247<=a_1;
mulc_2_247 : entity work.gfmul
port map(
a=>a_2,
b=>"111111010",
X=>mulr_2_247);

mulr_1_248<=a_1;
mulc_2_248 : entity work.gfmul
port map(
a=>a_2,
b=>"111100101",
X=>mulr_2_248);

mulr_1_249<=a_1;
mulc_2_249 : entity work.gfmul
port map(
a=>a_2,
b=>"111011011",
X=>mulr_2_249);

mulr_1_250<=a_1;
mulc_2_250 : entity work.gfmul
port map(
a=>a_2,
b=>"110100111",
X=>mulr_2_250);

mulr_1_251<=a_1;
mulc_2_251 : entity work.gfmul
port map(
a=>a_2,
b=>"101011111",
X=>mulr_2_251);

mulr_1_252<=a_1;
mulc_2_252 : entity work.gfmul
port map(
a=>a_2,
b=>"010101111",
X=>mulr_2_252);

mulr_1_253<=a_1;
mulc_2_253 : entity work.gfmul
port map(
a=>a_2,
b=>"101011110",
X=>mulr_2_253);

mulr_1_254<=a_1;
mulc_2_254 : entity work.gfmul
port map(
a=>a_2,
b=>"010101101",
X=>mulr_2_254);

mulr_1_255<=a_1;
mulc_2_255 : entity work.gfmul
port map(
a=>a_2,
b=>"101011010",
X=>mulr_2_255);

mulr_1_256<=a_1;
mulc_2_256 : entity work.gfmul
port map(
a=>a_2,
b=>"010100101",
X=>mulr_2_256);

mulr_1_257<=a_1;
mulc_2_257 : entity work.gfmul
port map(
a=>a_2,
b=>"101001010",
X=>mulr_2_257);

mulr_1_258<=a_1;
mulc_2_258 : entity work.gfmul
port map(
a=>a_2,
b=>"010000101",
X=>mulr_2_258);

mulr_1_259<=a_1;
mulc_2_259 : entity work.gfmul
port map(
a=>a_2,
b=>"100001010",
X=>mulr_2_259);

mulr_1_260<=a_1;
mulc_2_260 : entity work.gfmul
port map(
a=>a_2,
b=>"000000101",
X=>mulr_2_260);

mulr_1_261<=a_1;
mulc_2_261 : entity work.gfmul
port map(
a=>a_2,
b=>"000001010",
X=>mulr_2_261);

mulr_1_262<=a_1;
mulc_2_262 : entity work.gfmul
port map(
a=>a_2,
b=>"000010100",
X=>mulr_2_262);

mulr_1_263<=a_1;
mulc_2_263 : entity work.gfmul
port map(
a=>a_2,
b=>"000101000",
X=>mulr_2_263);

mulr_1_264<=a_1;
mulc_2_264 : entity work.gfmul
port map(
a=>a_2,
b=>"001010000",
X=>mulr_2_264);

mulr_1_265<=a_1;
mulc_2_265 : entity work.gfmul
port map(
a=>a_2,
b=>"010100000",
X=>mulr_2_265);

mulr_1_266<=a_1;
mulc_2_266 : entity work.gfmul
port map(
a=>a_2,
b=>"101000000",
X=>mulr_2_266);

mulr_1_267<=a_1;
mulc_2_267 : entity work.gfmul
port map(
a=>a_2,
b=>"010010001",
X=>mulr_2_267);

mulr_1_268<=a_1;
mulc_2_268 : entity work.gfmul
port map(
a=>a_2,
b=>"100100010",
X=>mulr_2_268);

mulr_1_269<=a_1;
mulc_2_269 : entity work.gfmul
port map(
a=>a_2,
b=>"001010101",
X=>mulr_2_269);

mulr_1_270<=a_1;
mulc_2_270 : entity work.gfmul
port map(
a=>a_2,
b=>"010101010",
X=>mulr_2_270);

mulr_1_271<=a_1;
mulc_2_271 : entity work.gfmul
port map(
a=>a_2,
b=>"101010100",
X=>mulr_2_271);

mulr_1_272<=a_1;
mulc_2_272 : entity work.gfmul
port map(
a=>a_2,
b=>"010111001",
X=>mulr_2_272);

mulr_1_273<=a_1;
mulc_2_273 : entity work.gfmul
port map(
a=>a_2,
b=>"101110010",
X=>mulr_2_273);

mulr_1_274<=a_1;
mulc_2_274 : entity work.gfmul
port map(
a=>a_2,
b=>"011110101",
X=>mulr_2_274);

mulr_1_275<=a_1;
mulc_2_275 : entity work.gfmul
port map(
a=>a_2,
b=>"111101010",
X=>mulr_2_275);

mulr_1_276<=a_1;
mulc_2_276 : entity work.gfmul
port map(
a=>a_2,
b=>"111000101",
X=>mulr_2_276);

mulr_1_277<=a_1;
mulc_2_277 : entity work.gfmul
port map(
a=>a_2,
b=>"110011011",
X=>mulr_2_277);

mulr_1_278<=a_1;
mulc_2_278 : entity work.gfmul
port map(
a=>a_2,
b=>"100100111",
X=>mulr_2_278);

mulr_1_279<=a_1;
mulc_2_279 : entity work.gfmul
port map(
a=>a_2,
b=>"001011111",
X=>mulr_2_279);

mulr_1_280<=a_1;
mulc_2_280 : entity work.gfmul
port map(
a=>a_2,
b=>"010111110",
X=>mulr_2_280);

mulr_1_281<=a_1;
mulc_2_281 : entity work.gfmul
port map(
a=>a_2,
b=>"101111100",
X=>mulr_2_281);

mulr_1_282<=a_1;
mulc_2_282 : entity work.gfmul
port map(
a=>a_2,
b=>"011101001",
X=>mulr_2_282);

mulr_1_283<=a_1;
mulc_2_283 : entity work.gfmul
port map(
a=>a_2,
b=>"111010010",
X=>mulr_2_283);

mulr_1_284<=a_1;
mulc_2_284 : entity work.gfmul
port map(
a=>a_2,
b=>"110110101",
X=>mulr_2_284);

mulr_1_285<=a_1;
mulc_2_285 : entity work.gfmul
port map(
a=>a_2,
b=>"101111011",
X=>mulr_2_285);

mulr_1_286<=a_1;
mulc_2_286 : entity work.gfmul
port map(
a=>a_2,
b=>"011100111",
X=>mulr_2_286);

mulr_1_287<=a_1;
mulc_2_287 : entity work.gfmul
port map(
a=>a_2,
b=>"111001110",
X=>mulr_2_287);

mulr_1_288<=a_1;
mulc_2_288 : entity work.gfmul
port map(
a=>a_2,
b=>"110001101",
X=>mulr_2_288);

mulr_1_289<=a_1;
mulc_2_289 : entity work.gfmul
port map(
a=>a_2,
b=>"100001011",
X=>mulr_2_289);

mulr_1_290<=a_1;
mulc_2_290 : entity work.gfmul
port map(
a=>a_2,
b=>"000000111",
X=>mulr_2_290);

mulr_1_291<=a_1;
mulc_2_291 : entity work.gfmul
port map(
a=>a_2,
b=>"000001110",
X=>mulr_2_291);

mulr_1_292<=a_1;
mulc_2_292 : entity work.gfmul
port map(
a=>a_2,
b=>"000011100",
X=>mulr_2_292);

mulr_1_293<=a_1;
mulc_2_293 : entity work.gfmul
port map(
a=>a_2,
b=>"000111000",
X=>mulr_2_293);

mulr_1_294<=a_1;
mulc_2_294 : entity work.gfmul
port map(
a=>a_2,
b=>"001110000",
X=>mulr_2_294);

mulr_1_295<=a_1;
mulc_2_295 : entity work.gfmul
port map(
a=>a_2,
b=>"011100000",
X=>mulr_2_295);

mulr_1_296<=a_1;
mulc_2_296 : entity work.gfmul
port map(
a=>a_2,
b=>"111000000",
X=>mulr_2_296);

mulr_1_297<=a_1;
mulc_2_297 : entity work.gfmul
port map(
a=>a_2,
b=>"110010001",
X=>mulr_2_297);

mulr_1_298<=a_1;
mulc_2_298 : entity work.gfmul
port map(
a=>a_2,
b=>"100110011",
X=>mulr_2_298);

mulr_1_299<=a_1;
mulc_2_299 : entity work.gfmul
port map(
a=>a_2,
b=>"001110111",
X=>mulr_2_299);

mulr_1_300<=a_1;
mulc_2_300 : entity work.gfmul
port map(
a=>a_2,
b=>"011101110",
X=>mulr_2_300);

mulr_1_301<=a_1;
mulc_2_301 : entity work.gfmul
port map(
a=>a_2,
b=>"111011100",
X=>mulr_2_301);

mulr_1_302<=a_1;
mulc_2_302 : entity work.gfmul
port map(
a=>a_2,
b=>"110101001",
X=>mulr_2_302);

mulr_1_303<=a_1;
mulc_2_303 : entity work.gfmul
port map(
a=>a_2,
b=>"101000011",
X=>mulr_2_303);

mulr_1_304<=a_1;
mulc_2_304 : entity work.gfmul
port map(
a=>a_2,
b=>"010010111",
X=>mulr_2_304);

mulr_1_305<=a_1;
mulc_2_305 : entity work.gfmul
port map(
a=>a_2,
b=>"100101110",
X=>mulr_2_305);

mulr_1_306<=a_1;
mulc_2_306 : entity work.gfmul
port map(
a=>a_2,
b=>"001001101",
X=>mulr_2_306);

mulr_1_307<=a_1;
mulc_2_307 : entity work.gfmul
port map(
a=>a_2,
b=>"010011010",
X=>mulr_2_307);

mulr_1_308<=a_1;
mulc_2_308 : entity work.gfmul
port map(
a=>a_2,
b=>"100110100",
X=>mulr_2_308);

mulr_1_309<=a_1;
mulc_2_309 : entity work.gfmul
port map(
a=>a_2,
b=>"001111001",
X=>mulr_2_309);

mulr_1_310<=a_1;
mulc_2_310 : entity work.gfmul
port map(
a=>a_2,
b=>"011110010",
X=>mulr_2_310);

mulr_1_311<=a_1;
mulc_2_311 : entity work.gfmul
port map(
a=>a_2,
b=>"111100100",
X=>mulr_2_311);

mulr_1_312<=a_1;
mulc_2_312 : entity work.gfmul
port map(
a=>a_2,
b=>"111011001",
X=>mulr_2_312);

mulr_1_313<=a_1;
mulc_2_313 : entity work.gfmul
port map(
a=>a_2,
b=>"110100011",
X=>mulr_2_313);

mulr_1_314<=a_1;
mulc_2_314 : entity work.gfmul
port map(
a=>a_2,
b=>"101010111",
X=>mulr_2_314);

mulr_1_315<=a_1;
mulc_2_315 : entity work.gfmul
port map(
a=>a_2,
b=>"010111111",
X=>mulr_2_315);

mulr_1_316<=a_1;
mulc_2_316 : entity work.gfmul
port map(
a=>a_2,
b=>"101111110",
X=>mulr_2_316);

mulr_1_317<=a_1;
mulc_2_317 : entity work.gfmul
port map(
a=>a_2,
b=>"011101101",
X=>mulr_2_317);

mulr_1_318<=a_1;
mulc_2_318 : entity work.gfmul
port map(
a=>a_2,
b=>"111011010",
X=>mulr_2_318);

mulr_1_319<=a_1;
mulc_2_319 : entity work.gfmul
port map(
a=>a_2,
b=>"110100101",
X=>mulr_2_319);

mulr_1_320<=a_1;
mulc_2_320 : entity work.gfmul
port map(
a=>a_2,
b=>"101011011",
X=>mulr_2_320);

mulr_1_321<=a_1;
mulc_2_321 : entity work.gfmul
port map(
a=>a_2,
b=>"010100111",
X=>mulr_2_321);

mulr_1_322<=a_1;
mulc_2_322 : entity work.gfmul
port map(
a=>a_2,
b=>"101001110",
X=>mulr_2_322);

mulr_1_323<=a_1;
mulc_2_323 : entity work.gfmul
port map(
a=>a_2,
b=>"010001101",
X=>mulr_2_323);

mulr_1_324<=a_1;
mulc_2_324 : entity work.gfmul
port map(
a=>a_2,
b=>"100011010",
X=>mulr_2_324);

mulr_1_325<=a_1;
mulc_2_325 : entity work.gfmul
port map(
a=>a_2,
b=>"000100101",
X=>mulr_2_325);

mulr_1_326<=a_1;
mulc_2_326 : entity work.gfmul
port map(
a=>a_2,
b=>"001001010",
X=>mulr_2_326);

mulr_1_327<=a_1;
mulc_2_327 : entity work.gfmul
port map(
a=>a_2,
b=>"010010100",
X=>mulr_2_327);

mulr_1_328<=a_1;
mulc_2_328 : entity work.gfmul
port map(
a=>a_2,
b=>"100101000",
X=>mulr_2_328);

mulr_1_329<=a_1;
mulc_2_329 : entity work.gfmul
port map(
a=>a_2,
b=>"001000001",
X=>mulr_2_329);

mulr_1_330<=a_1;
mulc_2_330 : entity work.gfmul
port map(
a=>a_2,
b=>"010000010",
X=>mulr_2_330);

mulr_1_331<=a_1;
mulc_2_331 : entity work.gfmul
port map(
a=>a_2,
b=>"100000100",
X=>mulr_2_331);

mulr_1_332<=a_1;
mulc_2_332 : entity work.gfmul
port map(
a=>a_2,
b=>"000011001",
X=>mulr_2_332);

mulr_1_333<=a_1;
mulc_2_333 : entity work.gfmul
port map(
a=>a_2,
b=>"000110010",
X=>mulr_2_333);

mulr_1_334<=a_1;
mulc_2_334 : entity work.gfmul
port map(
a=>a_2,
b=>"001100100",
X=>mulr_2_334);

mulr_1_335<=a_1;
mulc_2_335 : entity work.gfmul
port map(
a=>a_2,
b=>"011001000",
X=>mulr_2_335);

mulr_1_336<=a_1;
mulc_2_336 : entity work.gfmul
port map(
a=>a_2,
b=>"110010000",
X=>mulr_2_336);

mulr_1_337<=a_1;
mulc_2_337 : entity work.gfmul
port map(
a=>a_2,
b=>"100110001",
X=>mulr_2_337);

mulr_1_338<=a_1;
mulc_2_338 : entity work.gfmul
port map(
a=>a_2,
b=>"001110011",
X=>mulr_2_338);

mulr_1_339<=a_1;
mulc_2_339 : entity work.gfmul
port map(
a=>a_2,
b=>"011100110",
X=>mulr_2_339);

mulr_1_340<=a_1;
mulc_2_340 : entity work.gfmul
port map(
a=>a_2,
b=>"111001100",
X=>mulr_2_340);

mulr_1_341<=a_1;
mulc_2_341 : entity work.gfmul
port map(
a=>a_2,
b=>"110001001",
X=>mulr_2_341);

mulr_1_342<=a_1;
mulc_2_342 : entity work.gfmul
port map(
a=>a_2,
b=>"100000011",
X=>mulr_2_342);

mulr_1_343<=a_1;
mulc_2_343 : entity work.gfmul
port map(
a=>a_2,
b=>"000010111",
X=>mulr_2_343);

mulr_1_344<=a_1;
mulc_2_344 : entity work.gfmul
port map(
a=>a_2,
b=>"000101110",
X=>mulr_2_344);

mulr_1_345<=a_1;
mulc_2_345 : entity work.gfmul
port map(
a=>a_2,
b=>"001011100",
X=>mulr_2_345);

mulr_1_346<=a_1;
mulc_2_346 : entity work.gfmul
port map(
a=>a_2,
b=>"010111000",
X=>mulr_2_346);

mulr_1_347<=a_1;
mulc_2_347 : entity work.gfmul
port map(
a=>a_2,
b=>"101110000",
X=>mulr_2_347);

mulr_1_348<=a_1;
mulc_2_348 : entity work.gfmul
port map(
a=>a_2,
b=>"011110001",
X=>mulr_2_348);

mulr_1_349<=a_1;
mulc_2_349 : entity work.gfmul
port map(
a=>a_2,
b=>"111100010",
X=>mulr_2_349);

mulr_1_350<=a_1;
mulc_2_350 : entity work.gfmul
port map(
a=>a_2,
b=>"111010101",
X=>mulr_2_350);

mulr_1_351<=a_1;
mulc_2_351 : entity work.gfmul
port map(
a=>a_2,
b=>"110111011",
X=>mulr_2_351);

mulr_1_352<=a_1;
mulc_2_352 : entity work.gfmul
port map(
a=>a_2,
b=>"101100111",
X=>mulr_2_352);

mulr_1_353<=a_1;
mulc_2_353 : entity work.gfmul
port map(
a=>a_2,
b=>"011011111",
X=>mulr_2_353);

mulr_1_354<=a_1;
mulc_2_354 : entity work.gfmul
port map(
a=>a_2,
b=>"110111110",
X=>mulr_2_354);

mulr_1_355<=a_1;
mulc_2_355 : entity work.gfmul
port map(
a=>a_2,
b=>"101101101",
X=>mulr_2_355);

mulr_1_356<=a_1;
mulc_2_356 : entity work.gfmul
port map(
a=>a_2,
b=>"011001011",
X=>mulr_2_356);

mulr_1_357<=a_1;
mulc_2_357 : entity work.gfmul
port map(
a=>a_2,
b=>"110010110",
X=>mulr_2_357);

mulr_1_358<=a_1;
mulc_2_358 : entity work.gfmul
port map(
a=>a_2,
b=>"100111101",
X=>mulr_2_358);

mulr_1_359<=a_1;
mulc_2_359 : entity work.gfmul
port map(
a=>a_2,
b=>"001101011",
X=>mulr_2_359);

mulr_1_360<=a_1;
mulc_2_360 : entity work.gfmul
port map(
a=>a_2,
b=>"011010110",
X=>mulr_2_360);

mulr_1_361<=a_1;
mulc_2_361 : entity work.gfmul
port map(
a=>a_2,
b=>"110101100",
X=>mulr_2_361);

mulr_1_362<=a_1;
mulc_2_362 : entity work.gfmul
port map(
a=>a_2,
b=>"101001001",
X=>mulr_2_362);

mulr_1_363<=a_1;
mulc_2_363 : entity work.gfmul
port map(
a=>a_2,
b=>"010000011",
X=>mulr_2_363);

mulr_1_364<=a_1;
mulc_2_364 : entity work.gfmul
port map(
a=>a_2,
b=>"100000110",
X=>mulr_2_364);

mulr_1_365<=a_1;
mulc_2_365 : entity work.gfmul
port map(
a=>a_2,
b=>"000011101",
X=>mulr_2_365);

mulr_1_366<=a_1;
mulc_2_366 : entity work.gfmul
port map(
a=>a_2,
b=>"000111010",
X=>mulr_2_366);

mulr_1_367<=a_1;
mulc_2_367 : entity work.gfmul
port map(
a=>a_2,
b=>"001110100",
X=>mulr_2_367);

mulr_1_368<=a_1;
mulc_2_368 : entity work.gfmul
port map(
a=>a_2,
b=>"011101000",
X=>mulr_2_368);

mulr_1_369<=a_1;
mulc_2_369 : entity work.gfmul
port map(
a=>a_2,
b=>"111010000",
X=>mulr_2_369);

mulr_1_370<=a_1;
mulc_2_370 : entity work.gfmul
port map(
a=>a_2,
b=>"110110001",
X=>mulr_2_370);

mulr_1_371<=a_1;
mulc_2_371 : entity work.gfmul
port map(
a=>a_2,
b=>"101110011",
X=>mulr_2_371);

mulr_1_372<=a_1;
mulc_2_372 : entity work.gfmul
port map(
a=>a_2,
b=>"011110111",
X=>mulr_2_372);

mulr_1_373<=a_1;
mulc_2_373 : entity work.gfmul
port map(
a=>a_2,
b=>"111101110",
X=>mulr_2_373);

mulr_1_374<=a_1;
mulc_2_374 : entity work.gfmul
port map(
a=>a_2,
b=>"111001101",
X=>mulr_2_374);

mulr_1_375<=a_1;
mulc_2_375 : entity work.gfmul
port map(
a=>a_2,
b=>"110001011",
X=>mulr_2_375);

mulr_1_376<=a_1;
mulc_2_376 : entity work.gfmul
port map(
a=>a_2,
b=>"100000111",
X=>mulr_2_376);

mulr_1_377<=a_1;
mulc_2_377 : entity work.gfmul
port map(
a=>a_2,
b=>"000011111",
X=>mulr_2_377);

mulr_1_378<=a_1;
mulc_2_378 : entity work.gfmul
port map(
a=>a_2,
b=>"000111110",
X=>mulr_2_378);

mulr_1_379<=a_1;
mulc_2_379 : entity work.gfmul
port map(
a=>a_2,
b=>"001111100",
X=>mulr_2_379);

mulr_1_380<=a_1;
mulc_2_380 : entity work.gfmul
port map(
a=>a_2,
b=>"011111000",
X=>mulr_2_380);

mulr_1_381<=a_1;
mulc_2_381 : entity work.gfmul
port map(
a=>a_2,
b=>"111110000",
X=>mulr_2_381);

mulr_1_382<=a_1;
mulc_2_382 : entity work.gfmul
port map(
a=>a_2,
b=>"111110001",
X=>mulr_2_382);

mulr_1_383<=a_1;
mulc_2_383 : entity work.gfmul
port map(
a=>a_2,
b=>"111110011",
X=>mulr_2_383);

mulr_1_384<=a_1;
mulc_2_384 : entity work.gfmul
port map(
a=>a_2,
b=>"111110111",
X=>mulr_2_384);

mulr_1_385<=a_1;
mulc_2_385 : entity work.gfmul
port map(
a=>a_2,
b=>"111111111",
X=>mulr_2_385);

mulr_1_386<=a_1;
mulc_2_386 : entity work.gfmul
port map(
a=>a_2,
b=>"111101111",
X=>mulr_2_386);

mulr_1_387<=a_1;
mulc_2_387 : entity work.gfmul
port map(
a=>a_2,
b=>"111001111",
X=>mulr_2_387);

mulr_1_388<=a_1;
mulc_2_388 : entity work.gfmul
port map(
a=>a_2,
b=>"110001111",
X=>mulr_2_388);

mulr_1_389<=a_1;
mulc_2_389 : entity work.gfmul
port map(
a=>a_2,
b=>"100001111",
X=>mulr_2_389);

mulr_1_390<=a_1;
mulc_2_390 : entity work.gfmul
port map(
a=>a_2,
b=>"000001111",
X=>mulr_2_390);

mulr_1_391<=a_1;
mulc_2_391 : entity work.gfmul
port map(
a=>a_2,
b=>"000011110",
X=>mulr_2_391);

mulr_1_392<=a_1;
mulc_2_392 : entity work.gfmul
port map(
a=>a_2,
b=>"000111100",
X=>mulr_2_392);

mulr_1_393<=a_1;
mulc_2_393 : entity work.gfmul
port map(
a=>a_2,
b=>"001111000",
X=>mulr_2_393);

mulr_1_394<=a_1;
mulc_2_394 : entity work.gfmul
port map(
a=>a_2,
b=>"011110000",
X=>mulr_2_394);

mulr_1_395<=a_1;
mulc_2_395 : entity work.gfmul
port map(
a=>a_2,
b=>"111100000",
X=>mulr_2_395);

mulr_1_396<=a_1;
mulc_2_396 : entity work.gfmul
port map(
a=>a_2,
b=>"111010001",
X=>mulr_2_396);

mulr_1_397<=a_1;
mulc_2_397 : entity work.gfmul
port map(
a=>a_2,
b=>"110110011",
X=>mulr_2_397);

mulr_1_398<=a_1;
mulc_2_398 : entity work.gfmul
port map(
a=>a_2,
b=>"101110111",
X=>mulr_2_398);

mulr_1_399<=a_1;
mulc_2_399 : entity work.gfmul
port map(
a=>a_2,
b=>"011111111",
X=>mulr_2_399);

mulr_1_400<=a_1;
mulc_2_400 : entity work.gfmul
port map(
a=>a_2,
b=>"111111110",
X=>mulr_2_400);

mulr_1_401<=a_1;
mulc_2_401 : entity work.gfmul
port map(
a=>a_2,
b=>"111101101",
X=>mulr_2_401);

mulr_1_402<=a_1;
mulc_2_402 : entity work.gfmul
port map(
a=>a_2,
b=>"111001011",
X=>mulr_2_402);

mulr_1_403<=a_1;
mulc_2_403 : entity work.gfmul
port map(
a=>a_2,
b=>"110000111",
X=>mulr_2_403);

mulr_1_404<=a_1;
mulc_2_404 : entity work.gfmul
port map(
a=>a_2,
b=>"100011111",
X=>mulr_2_404);

mulr_1_405<=a_1;
mulc_2_405 : entity work.gfmul
port map(
a=>a_2,
b=>"000101111",
X=>mulr_2_405);

mulr_1_406<=a_1;
mulc_2_406 : entity work.gfmul
port map(
a=>a_2,
b=>"001011110",
X=>mulr_2_406);

mulr_1_407<=a_1;
mulc_2_407 : entity work.gfmul
port map(
a=>a_2,
b=>"010111100",
X=>mulr_2_407);

mulr_1_408<=a_1;
mulc_2_408 : entity work.gfmul
port map(
a=>a_2,
b=>"101111000",
X=>mulr_2_408);

mulr_1_409<=a_1;
mulc_2_409 : entity work.gfmul
port map(
a=>a_2,
b=>"011100001",
X=>mulr_2_409);

mulr_1_410<=a_1;
mulc_2_410 : entity work.gfmul
port map(
a=>a_2,
b=>"111000010",
X=>mulr_2_410);

mulr_1_411<=a_1;
mulc_2_411 : entity work.gfmul
port map(
a=>a_2,
b=>"110010101",
X=>mulr_2_411);

mulr_1_412<=a_1;
mulc_2_412 : entity work.gfmul
port map(
a=>a_2,
b=>"100111011",
X=>mulr_2_412);

mulr_1_413<=a_1;
mulc_2_413 : entity work.gfmul
port map(
a=>a_2,
b=>"001100111",
X=>mulr_2_413);

mulr_1_414<=a_1;
mulc_2_414 : entity work.gfmul
port map(
a=>a_2,
b=>"011001110",
X=>mulr_2_414);

mulr_1_415<=a_1;
mulc_2_415 : entity work.gfmul
port map(
a=>a_2,
b=>"110011100",
X=>mulr_2_415);

mulr_1_416<=a_1;
mulc_2_416 : entity work.gfmul
port map(
a=>a_2,
b=>"100101001",
X=>mulr_2_416);

mulr_1_417<=a_1;
mulc_2_417 : entity work.gfmul
port map(
a=>a_2,
b=>"001000011",
X=>mulr_2_417);

mulr_1_418<=a_1;
mulc_2_418 : entity work.gfmul
port map(
a=>a_2,
b=>"010000110",
X=>mulr_2_418);

mulr_1_419<=a_1;
mulc_2_419 : entity work.gfmul
port map(
a=>a_2,
b=>"100001100",
X=>mulr_2_419);

mulr_1_420<=a_1;
mulc_2_420 : entity work.gfmul
port map(
a=>a_2,
b=>"000001001",
X=>mulr_2_420);

mulr_1_421<=a_1;
mulc_2_421 : entity work.gfmul
port map(
a=>a_2,
b=>"000010010",
X=>mulr_2_421);

mulr_1_422<=a_1;
mulc_2_422 : entity work.gfmul
port map(
a=>a_2,
b=>"000100100",
X=>mulr_2_422);

mulr_1_423<=a_1;
mulc_2_423 : entity work.gfmul
port map(
a=>a_2,
b=>"001001000",
X=>mulr_2_423);

mulr_1_424<=a_1;
mulc_2_424 : entity work.gfmul
port map(
a=>a_2,
b=>"010010000",
X=>mulr_2_424);

mulr_1_425<=a_1;
mulc_2_425 : entity work.gfmul
port map(
a=>a_2,
b=>"100100000",
X=>mulr_2_425);

mulr_1_426<=a_1;
mulc_2_426 : entity work.gfmul
port map(
a=>a_2,
b=>"001010001",
X=>mulr_2_426);

mulr_1_427<=a_1;
mulc_2_427 : entity work.gfmul
port map(
a=>a_2,
b=>"010100010",
X=>mulr_2_427);

mulr_1_428<=a_1;
mulc_2_428 : entity work.gfmul
port map(
a=>a_2,
b=>"101000100",
X=>mulr_2_428);

mulr_1_429<=a_1;
mulc_2_429 : entity work.gfmul
port map(
a=>a_2,
b=>"010011001",
X=>mulr_2_429);

mulr_1_430<=a_1;
mulc_2_430 : entity work.gfmul
port map(
a=>a_2,
b=>"100110010",
X=>mulr_2_430);

mulr_1_431<=a_1;
mulc_2_431 : entity work.gfmul
port map(
a=>a_2,
b=>"001110101",
X=>mulr_2_431);

mulr_1_432<=a_1;
mulc_2_432 : entity work.gfmul
port map(
a=>a_2,
b=>"011101010",
X=>mulr_2_432);

mulr_1_433<=a_1;
mulc_2_433 : entity work.gfmul
port map(
a=>a_2,
b=>"111010100",
X=>mulr_2_433);

mulr_1_434<=a_1;
mulc_2_434 : entity work.gfmul
port map(
a=>a_2,
b=>"110111001",
X=>mulr_2_434);

mulr_1_435<=a_1;
mulc_2_435 : entity work.gfmul
port map(
a=>a_2,
b=>"101100011",
X=>mulr_2_435);

mulr_1_436<=a_1;
mulc_2_436 : entity work.gfmul
port map(
a=>a_2,
b=>"011010111",
X=>mulr_2_436);

mulr_1_437<=a_1;
mulc_2_437 : entity work.gfmul
port map(
a=>a_2,
b=>"110101110",
X=>mulr_2_437);

mulr_1_438<=a_1;
mulc_2_438 : entity work.gfmul
port map(
a=>a_2,
b=>"101001101",
X=>mulr_2_438);

mulr_1_439<=a_1;
mulc_2_439 : entity work.gfmul
port map(
a=>a_2,
b=>"010001011",
X=>mulr_2_439);

mulr_1_440<=a_1;
mulc_2_440 : entity work.gfmul
port map(
a=>a_2,
b=>"100010110",
X=>mulr_2_440);

mulr_1_441<=a_1;
mulc_2_441 : entity work.gfmul
port map(
a=>a_2,
b=>"000111101",
X=>mulr_2_441);

mulr_1_442<=a_1;
mulc_2_442 : entity work.gfmul
port map(
a=>a_2,
b=>"001111010",
X=>mulr_2_442);

mulr_1_443<=a_1;
mulc_2_443 : entity work.gfmul
port map(
a=>a_2,
b=>"011110100",
X=>mulr_2_443);

mulr_1_444<=a_1;
mulc_2_444 : entity work.gfmul
port map(
a=>a_2,
b=>"111101000",
X=>mulr_2_444);

mulr_1_445<=a_1;
mulc_2_445 : entity work.gfmul
port map(
a=>a_2,
b=>"111000001",
X=>mulr_2_445);

mulr_1_446<=a_1;
mulc_2_446 : entity work.gfmul
port map(
a=>a_2,
b=>"110010011",
X=>mulr_2_446);

mulr_1_447<=a_1;
mulc_2_447 : entity work.gfmul
port map(
a=>a_2,
b=>"100110111",
X=>mulr_2_447);

mulr_1_448<=a_1;
mulc_2_448 : entity work.gfmul
port map(
a=>a_2,
b=>"001111111",
X=>mulr_2_448);

mulr_1_449<=a_1;
mulc_2_449 : entity work.gfmul
port map(
a=>a_2,
b=>"011111110",
X=>mulr_2_449);

mulr_1_450<=a_1;
mulc_2_450 : entity work.gfmul
port map(
a=>a_2,
b=>"111111100",
X=>mulr_2_450);

mulr_1_451<=a_1;
mulc_2_451 : entity work.gfmul
port map(
a=>a_2,
b=>"111101001",
X=>mulr_2_451);

mulr_1_452<=a_1;
mulc_2_452 : entity work.gfmul
port map(
a=>a_2,
b=>"111000011",
X=>mulr_2_452);

mulr_1_453<=a_1;
mulc_2_453 : entity work.gfmul
port map(
a=>a_2,
b=>"110010111",
X=>mulr_2_453);

mulr_1_454<=a_1;
mulc_2_454 : entity work.gfmul
port map(
a=>a_2,
b=>"100111111",
X=>mulr_2_454);

mulr_1_455<=a_1;
mulc_2_455 : entity work.gfmul
port map(
a=>a_2,
b=>"001101111",
X=>mulr_2_455);

mulr_1_456<=a_1;
mulc_2_456 : entity work.gfmul
port map(
a=>a_2,
b=>"011011110",
X=>mulr_2_456);

mulr_1_457<=a_1;
mulc_2_457 : entity work.gfmul
port map(
a=>a_2,
b=>"110111100",
X=>mulr_2_457);

mulr_1_458<=a_1;
mulc_2_458 : entity work.gfmul
port map(
a=>a_2,
b=>"101101001",
X=>mulr_2_458);

mulr_1_459<=a_1;
mulc_2_459 : entity work.gfmul
port map(
a=>a_2,
b=>"011000011",
X=>mulr_2_459);

mulr_1_460<=a_1;
mulc_2_460 : entity work.gfmul
port map(
a=>a_2,
b=>"110000110",
X=>mulr_2_460);

mulr_1_461<=a_1;
mulc_2_461 : entity work.gfmul
port map(
a=>a_2,
b=>"100011101",
X=>mulr_2_461);

mulr_1_462<=a_1;
mulc_2_462 : entity work.gfmul
port map(
a=>a_2,
b=>"000101011",
X=>mulr_2_462);

mulr_1_463<=a_1;
mulc_2_463 : entity work.gfmul
port map(
a=>a_2,
b=>"001010110",
X=>mulr_2_463);

mulr_1_464<=a_1;
mulc_2_464 : entity work.gfmul
port map(
a=>a_2,
b=>"010101100",
X=>mulr_2_464);

mulr_1_465<=a_1;
mulc_2_465 : entity work.gfmul
port map(
a=>a_2,
b=>"101011000",
X=>mulr_2_465);

mulr_1_466<=a_1;
mulc_2_466 : entity work.gfmul
port map(
a=>a_2,
b=>"010100001",
X=>mulr_2_466);

mulr_1_467<=a_1;
mulc_2_467 : entity work.gfmul
port map(
a=>a_2,
b=>"101000010",
X=>mulr_2_467);

mulr_1_468<=a_1;
mulc_2_468 : entity work.gfmul
port map(
a=>a_2,
b=>"010010101",
X=>mulr_2_468);

mulr_1_469<=a_1;
mulc_2_469 : entity work.gfmul
port map(
a=>a_2,
b=>"100101010",
X=>mulr_2_469);

mulr_1_470<=a_1;
mulc_2_470 : entity work.gfmul
port map(
a=>a_2,
b=>"001000101",
X=>mulr_2_470);

mulr_1_471<=a_1;
mulc_2_471 : entity work.gfmul
port map(
a=>a_2,
b=>"010001010",
X=>mulr_2_471);

mulr_1_472<=a_1;
mulc_2_472 : entity work.gfmul
port map(
a=>a_2,
b=>"100010100",
X=>mulr_2_472);

mulr_1_473<=a_1;
mulc_2_473 : entity work.gfmul
port map(
a=>a_2,
b=>"000111001",
X=>mulr_2_473);

mulr_1_474<=a_1;
mulc_2_474 : entity work.gfmul
port map(
a=>a_2,
b=>"001110010",
X=>mulr_2_474);

mulr_1_475<=a_1;
mulc_2_475 : entity work.gfmul
port map(
a=>a_2,
b=>"011100100",
X=>mulr_2_475);

mulr_1_476<=a_1;
mulc_2_476 : entity work.gfmul
port map(
a=>a_2,
b=>"111001000",
X=>mulr_2_476);

mulr_1_477<=a_1;
mulc_2_477 : entity work.gfmul
port map(
a=>a_2,
b=>"110000001",
X=>mulr_2_477);

mulr_1_478<=a_1;
mulc_2_478 : entity work.gfmul
port map(
a=>a_2,
b=>"100010011",
X=>mulr_2_478);

mulr_1_479<=a_1;
mulc_2_479 : entity work.gfmul
port map(
a=>a_2,
b=>"000110111",
X=>mulr_2_479);

mulr_1_480<=a_1;
mulc_2_480 : entity work.gfmul
port map(
a=>a_2,
b=>"001101110",
X=>mulr_2_480);

mulr_1_481<=a_1;
mulc_2_481 : entity work.gfmul
port map(
a=>a_2,
b=>"011011100",
X=>mulr_2_481);

mulr_1_482<=a_1;
mulc_2_482 : entity work.gfmul
port map(
a=>a_2,
b=>"110111000",
X=>mulr_2_482);

mulr_1_483<=a_1;
mulc_2_483 : entity work.gfmul
port map(
a=>a_2,
b=>"101100001",
X=>mulr_2_483);

mulr_1_484<=a_1;
mulc_2_484 : entity work.gfmul
port map(
a=>a_2,
b=>"011010011",
X=>mulr_2_484);

mulr_1_485<=a_1;
mulc_2_485 : entity work.gfmul
port map(
a=>a_2,
b=>"110100110",
X=>mulr_2_485);

mulr_1_486<=a_1;
mulc_2_486 : entity work.gfmul
port map(
a=>a_2,
b=>"101011101",
X=>mulr_2_486);

mulr_1_487<=a_1;
mulc_2_487 : entity work.gfmul
port map(
a=>a_2,
b=>"010101011",
X=>mulr_2_487);

mulr_1_488<=a_1;
mulc_2_488 : entity work.gfmul
port map(
a=>a_2,
b=>"101010110",
X=>mulr_2_488);

mulr_1_489<=a_1;
mulc_2_489 : entity work.gfmul
port map(
a=>a_2,
b=>"010111101",
X=>mulr_2_489);

mulr_1_490<=a_1;
mulc_2_490 : entity work.gfmul
port map(
a=>a_2,
b=>"101111010",
X=>mulr_2_490);

mulr_1_491<=a_1;
mulc_2_491 : entity work.gfmul
port map(
a=>a_2,
b=>"011100101",
X=>mulr_2_491);

mulr_1_492<=a_1;
mulc_2_492 : entity work.gfmul
port map(
a=>a_2,
b=>"111001010",
X=>mulr_2_492);

mulr_1_493<=a_1;
mulc_2_493 : entity work.gfmul
port map(
a=>a_2,
b=>"110000101",
X=>mulr_2_493);

mulr_1_494<=a_1;
mulc_2_494 : entity work.gfmul
port map(
a=>a_2,
b=>"100011011",
X=>mulr_2_494);

mulr_1_495<=a_1;
mulc_2_495 : entity work.gfmul
port map(
a=>a_2,
b=>"000100111",
X=>mulr_2_495);

mulr_1_496<=a_1;
mulc_2_496 : entity work.gfmul
port map(
a=>a_2,
b=>"001001110",
X=>mulr_2_496);

mulr_1_497<=a_1;
mulc_2_497 : entity work.gfmul
port map(
a=>a_2,
b=>"010011100",
X=>mulr_2_497);

mulr_1_498<=a_1;
mulc_2_498 : entity work.gfmul
port map(
a=>a_2,
b=>"100111000",
X=>mulr_2_498);

mulr_1_499<=a_1;
mulc_2_499 : entity work.gfmul
port map(
a=>a_2,
b=>"001100001",
X=>mulr_2_499);

mulr_1_500<=a_1;
mulc_2_500 : entity work.gfmul
port map(
a=>a_2,
b=>"011000010",
X=>mulr_2_500);

mulr_1_501<=a_1;
mulc_2_501 : entity work.gfmul
port map(
a=>a_2,
b=>"110000100",
X=>mulr_2_501);

mulr_1_502<=a_1;
mulc_2_502 : entity work.gfmul
port map(
a=>a_2,
b=>"100011001",
X=>mulr_2_502);

mulr_1_503<=a_1;
mulc_2_503 : entity work.gfmul
port map(
a=>a_2,
b=>"000100011",
X=>mulr_2_503);

mulr_1_504<=a_1;
mulc_2_504 : entity work.gfmul
port map(
a=>a_2,
b=>"001000110",
X=>mulr_2_504);

mulr_1_505<=a_1;
mulc_2_505 : entity work.gfmul
port map(
a=>a_2,
b=>"010001100",
X=>mulr_2_505);

mulr_1_506<=a_1;
mulc_2_506 : entity work.gfmul
port map(
a=>a_2,
b=>"100011000",
X=>mulr_2_506);

mulr_1_507<=a_1;
mulc_2_507 : entity work.gfmul
port map(
a=>a_2,
b=>"000100001",
X=>mulr_2_507);

mulr_1_508<=a_1;
mulc_2_508 : entity work.gfmul
port map(
a=>a_2,
b=>"001000010",
X=>mulr_2_508);

mulr_1_509<=a_1;
mulc_2_509 : entity work.gfmul
port map(
a=>a_2,
b=>"010000100",
X=>mulr_2_509);

mulr_1_510<=a_1;
mulc_2_510 : entity work.gfmul
port map(
a=>a_2,
b=>"100001000",
X=>mulr_2_510);

mulr_1_511<=a_1;
mulc_2_511 : entity work.gfmul
port map(
a=>a_2,
b=>"000000001",
X=>mulr_2_511);

sumr_1<= mulr_1_1 xor mulr_2_1;
sumr_2<= mulr_1_2 xor mulr_2_2;
sumr_3<= mulr_1_3 xor mulr_2_3;
sumr_4<= mulr_1_4 xor mulr_2_4;
sumr_5<= mulr_1_5 xor mulr_2_5;
sumr_6<= mulr_1_6 xor mulr_2_6;
sumr_7<= mulr_1_7 xor mulr_2_7;
sumr_8<= mulr_1_8 xor mulr_2_8;
sumr_9<= mulr_1_9 xor mulr_2_9;
sumr_10<= mulr_1_10 xor mulr_2_10;
sumr_11<= mulr_1_11 xor mulr_2_11;
sumr_12<= mulr_1_12 xor mulr_2_12;
sumr_13<= mulr_1_13 xor mulr_2_13;
sumr_14<= mulr_1_14 xor mulr_2_14;
sumr_15<= mulr_1_15 xor mulr_2_15;
sumr_16<= mulr_1_16 xor mulr_2_16;
sumr_17<= mulr_1_17 xor mulr_2_17;
sumr_18<= mulr_1_18 xor mulr_2_18;
sumr_19<= mulr_1_19 xor mulr_2_19;
sumr_20<= mulr_1_20 xor mulr_2_20;
sumr_21<= mulr_1_21 xor mulr_2_21;
sumr_22<= mulr_1_22 xor mulr_2_22;
sumr_23<= mulr_1_23 xor mulr_2_23;
sumr_24<= mulr_1_24 xor mulr_2_24;
sumr_25<= mulr_1_25 xor mulr_2_25;
sumr_26<= mulr_1_26 xor mulr_2_26;
sumr_27<= mulr_1_27 xor mulr_2_27;
sumr_28<= mulr_1_28 xor mulr_2_28;
sumr_29<= mulr_1_29 xor mulr_2_29;
sumr_30<= mulr_1_30 xor mulr_2_30;
sumr_31<= mulr_1_31 xor mulr_2_31;
sumr_32<= mulr_1_32 xor mulr_2_32;
sumr_33<= mulr_1_33 xor mulr_2_33;
sumr_34<= mulr_1_34 xor mulr_2_34;
sumr_35<= mulr_1_35 xor mulr_2_35;
sumr_36<= mulr_1_36 xor mulr_2_36;
sumr_37<= mulr_1_37 xor mulr_2_37;
sumr_38<= mulr_1_38 xor mulr_2_38;
sumr_39<= mulr_1_39 xor mulr_2_39;
sumr_40<= mulr_1_40 xor mulr_2_40;
sumr_41<= mulr_1_41 xor mulr_2_41;
sumr_42<= mulr_1_42 xor mulr_2_42;
sumr_43<= mulr_1_43 xor mulr_2_43;
sumr_44<= mulr_1_44 xor mulr_2_44;
sumr_45<= mulr_1_45 xor mulr_2_45;
sumr_46<= mulr_1_46 xor mulr_2_46;
sumr_47<= mulr_1_47 xor mulr_2_47;
sumr_48<= mulr_1_48 xor mulr_2_48;
sumr_49<= mulr_1_49 xor mulr_2_49;
sumr_50<= mulr_1_50 xor mulr_2_50;
sumr_51<= mulr_1_51 xor mulr_2_51;
sumr_52<= mulr_1_52 xor mulr_2_52;
sumr_53<= mulr_1_53 xor mulr_2_53;
sumr_54<= mulr_1_54 xor mulr_2_54;
sumr_55<= mulr_1_55 xor mulr_2_55;
sumr_56<= mulr_1_56 xor mulr_2_56;
sumr_57<= mulr_1_57 xor mulr_2_57;
sumr_58<= mulr_1_58 xor mulr_2_58;
sumr_59<= mulr_1_59 xor mulr_2_59;
sumr_60<= mulr_1_60 xor mulr_2_60;
sumr_61<= mulr_1_61 xor mulr_2_61;
sumr_62<= mulr_1_62 xor mulr_2_62;
sumr_63<= mulr_1_63 xor mulr_2_63;
sumr_64<= mulr_1_64 xor mulr_2_64;
sumr_65<= mulr_1_65 xor mulr_2_65;
sumr_66<= mulr_1_66 xor mulr_2_66;
sumr_67<= mulr_1_67 xor mulr_2_67;
sumr_68<= mulr_1_68 xor mulr_2_68;
sumr_69<= mulr_1_69 xor mulr_2_69;
sumr_70<= mulr_1_70 xor mulr_2_70;
sumr_71<= mulr_1_71 xor mulr_2_71;
sumr_72<= mulr_1_72 xor mulr_2_72;
sumr_73<= mulr_1_73 xor mulr_2_73;
sumr_74<= mulr_1_74 xor mulr_2_74;
sumr_75<= mulr_1_75 xor mulr_2_75;
sumr_76<= mulr_1_76 xor mulr_2_76;
sumr_77<= mulr_1_77 xor mulr_2_77;
sumr_78<= mulr_1_78 xor mulr_2_78;
sumr_79<= mulr_1_79 xor mulr_2_79;
sumr_80<= mulr_1_80 xor mulr_2_80;
sumr_81<= mulr_1_81 xor mulr_2_81;
sumr_82<= mulr_1_82 xor mulr_2_82;
sumr_83<= mulr_1_83 xor mulr_2_83;
sumr_84<= mulr_1_84 xor mulr_2_84;
sumr_85<= mulr_1_85 xor mulr_2_85;
sumr_86<= mulr_1_86 xor mulr_2_86;
sumr_87<= mulr_1_87 xor mulr_2_87;
sumr_88<= mulr_1_88 xor mulr_2_88;
sumr_89<= mulr_1_89 xor mulr_2_89;
sumr_90<= mulr_1_90 xor mulr_2_90;
sumr_91<= mulr_1_91 xor mulr_2_91;
sumr_92<= mulr_1_92 xor mulr_2_92;
sumr_93<= mulr_1_93 xor mulr_2_93;
sumr_94<= mulr_1_94 xor mulr_2_94;
sumr_95<= mulr_1_95 xor mulr_2_95;
sumr_96<= mulr_1_96 xor mulr_2_96;
sumr_97<= mulr_1_97 xor mulr_2_97;
sumr_98<= mulr_1_98 xor mulr_2_98;
sumr_99<= mulr_1_99 xor mulr_2_99;
sumr_100<= mulr_1_100 xor mulr_2_100;
sumr_101<= mulr_1_101 xor mulr_2_101;
sumr_102<= mulr_1_102 xor mulr_2_102;
sumr_103<= mulr_1_103 xor mulr_2_103;
sumr_104<= mulr_1_104 xor mulr_2_104;
sumr_105<= mulr_1_105 xor mulr_2_105;
sumr_106<= mulr_1_106 xor mulr_2_106;
sumr_107<= mulr_1_107 xor mulr_2_107;
sumr_108<= mulr_1_108 xor mulr_2_108;
sumr_109<= mulr_1_109 xor mulr_2_109;
sumr_110<= mulr_1_110 xor mulr_2_110;
sumr_111<= mulr_1_111 xor mulr_2_111;
sumr_112<= mulr_1_112 xor mulr_2_112;
sumr_113<= mulr_1_113 xor mulr_2_113;
sumr_114<= mulr_1_114 xor mulr_2_114;
sumr_115<= mulr_1_115 xor mulr_2_115;
sumr_116<= mulr_1_116 xor mulr_2_116;
sumr_117<= mulr_1_117 xor mulr_2_117;
sumr_118<= mulr_1_118 xor mulr_2_118;
sumr_119<= mulr_1_119 xor mulr_2_119;
sumr_120<= mulr_1_120 xor mulr_2_120;
sumr_121<= mulr_1_121 xor mulr_2_121;
sumr_122<= mulr_1_122 xor mulr_2_122;
sumr_123<= mulr_1_123 xor mulr_2_123;
sumr_124<= mulr_1_124 xor mulr_2_124;
sumr_125<= mulr_1_125 xor mulr_2_125;
sumr_126<= mulr_1_126 xor mulr_2_126;
sumr_127<= mulr_1_127 xor mulr_2_127;
sumr_128<= mulr_1_128 xor mulr_2_128;
sumr_129<= mulr_1_129 xor mulr_2_129;
sumr_130<= mulr_1_130 xor mulr_2_130;
sumr_131<= mulr_1_131 xor mulr_2_131;
sumr_132<= mulr_1_132 xor mulr_2_132;
sumr_133<= mulr_1_133 xor mulr_2_133;
sumr_134<= mulr_1_134 xor mulr_2_134;
sumr_135<= mulr_1_135 xor mulr_2_135;
sumr_136<= mulr_1_136 xor mulr_2_136;
sumr_137<= mulr_1_137 xor mulr_2_137;
sumr_138<= mulr_1_138 xor mulr_2_138;
sumr_139<= mulr_1_139 xor mulr_2_139;
sumr_140<= mulr_1_140 xor mulr_2_140;
sumr_141<= mulr_1_141 xor mulr_2_141;
sumr_142<= mulr_1_142 xor mulr_2_142;
sumr_143<= mulr_1_143 xor mulr_2_143;
sumr_144<= mulr_1_144 xor mulr_2_144;
sumr_145<= mulr_1_145 xor mulr_2_145;
sumr_146<= mulr_1_146 xor mulr_2_146;
sumr_147<= mulr_1_147 xor mulr_2_147;
sumr_148<= mulr_1_148 xor mulr_2_148;
sumr_149<= mulr_1_149 xor mulr_2_149;
sumr_150<= mulr_1_150 xor mulr_2_150;
sumr_151<= mulr_1_151 xor mulr_2_151;
sumr_152<= mulr_1_152 xor mulr_2_152;
sumr_153<= mulr_1_153 xor mulr_2_153;
sumr_154<= mulr_1_154 xor mulr_2_154;
sumr_155<= mulr_1_155 xor mulr_2_155;
sumr_156<= mulr_1_156 xor mulr_2_156;
sumr_157<= mulr_1_157 xor mulr_2_157;
sumr_158<= mulr_1_158 xor mulr_2_158;
sumr_159<= mulr_1_159 xor mulr_2_159;
sumr_160<= mulr_1_160 xor mulr_2_160;
sumr_161<= mulr_1_161 xor mulr_2_161;
sumr_162<= mulr_1_162 xor mulr_2_162;
sumr_163<= mulr_1_163 xor mulr_2_163;
sumr_164<= mulr_1_164 xor mulr_2_164;
sumr_165<= mulr_1_165 xor mulr_2_165;
sumr_166<= mulr_1_166 xor mulr_2_166;
sumr_167<= mulr_1_167 xor mulr_2_167;
sumr_168<= mulr_1_168 xor mulr_2_168;
sumr_169<= mulr_1_169 xor mulr_2_169;
sumr_170<= mulr_1_170 xor mulr_2_170;
sumr_171<= mulr_1_171 xor mulr_2_171;
sumr_172<= mulr_1_172 xor mulr_2_172;
sumr_173<= mulr_1_173 xor mulr_2_173;
sumr_174<= mulr_1_174 xor mulr_2_174;
sumr_175<= mulr_1_175 xor mulr_2_175;
sumr_176<= mulr_1_176 xor mulr_2_176;
sumr_177<= mulr_1_177 xor mulr_2_177;
sumr_178<= mulr_1_178 xor mulr_2_178;
sumr_179<= mulr_1_179 xor mulr_2_179;
sumr_180<= mulr_1_180 xor mulr_2_180;
sumr_181<= mulr_1_181 xor mulr_2_181;
sumr_182<= mulr_1_182 xor mulr_2_182;
sumr_183<= mulr_1_183 xor mulr_2_183;
sumr_184<= mulr_1_184 xor mulr_2_184;
sumr_185<= mulr_1_185 xor mulr_2_185;
sumr_186<= mulr_1_186 xor mulr_2_186;
sumr_187<= mulr_1_187 xor mulr_2_187;
sumr_188<= mulr_1_188 xor mulr_2_188;
sumr_189<= mulr_1_189 xor mulr_2_189;
sumr_190<= mulr_1_190 xor mulr_2_190;
sumr_191<= mulr_1_191 xor mulr_2_191;
sumr_192<= mulr_1_192 xor mulr_2_192;
sumr_193<= mulr_1_193 xor mulr_2_193;
sumr_194<= mulr_1_194 xor mulr_2_194;
sumr_195<= mulr_1_195 xor mulr_2_195;
sumr_196<= mulr_1_196 xor mulr_2_196;
sumr_197<= mulr_1_197 xor mulr_2_197;
sumr_198<= mulr_1_198 xor mulr_2_198;
sumr_199<= mulr_1_199 xor mulr_2_199;
sumr_200<= mulr_1_200 xor mulr_2_200;
sumr_201<= mulr_1_201 xor mulr_2_201;
sumr_202<= mulr_1_202 xor mulr_2_202;
sumr_203<= mulr_1_203 xor mulr_2_203;
sumr_204<= mulr_1_204 xor mulr_2_204;
sumr_205<= mulr_1_205 xor mulr_2_205;
sumr_206<= mulr_1_206 xor mulr_2_206;
sumr_207<= mulr_1_207 xor mulr_2_207;
sumr_208<= mulr_1_208 xor mulr_2_208;
sumr_209<= mulr_1_209 xor mulr_2_209;
sumr_210<= mulr_1_210 xor mulr_2_210;
sumr_211<= mulr_1_211 xor mulr_2_211;
sumr_212<= mulr_1_212 xor mulr_2_212;
sumr_213<= mulr_1_213 xor mulr_2_213;
sumr_214<= mulr_1_214 xor mulr_2_214;
sumr_215<= mulr_1_215 xor mulr_2_215;
sumr_216<= mulr_1_216 xor mulr_2_216;
sumr_217<= mulr_1_217 xor mulr_2_217;
sumr_218<= mulr_1_218 xor mulr_2_218;
sumr_219<= mulr_1_219 xor mulr_2_219;
sumr_220<= mulr_1_220 xor mulr_2_220;
sumr_221<= mulr_1_221 xor mulr_2_221;
sumr_222<= mulr_1_222 xor mulr_2_222;
sumr_223<= mulr_1_223 xor mulr_2_223;
sumr_224<= mulr_1_224 xor mulr_2_224;
sumr_225<= mulr_1_225 xor mulr_2_225;
sumr_226<= mulr_1_226 xor mulr_2_226;
sumr_227<= mulr_1_227 xor mulr_2_227;
sumr_228<= mulr_1_228 xor mulr_2_228;
sumr_229<= mulr_1_229 xor mulr_2_229;
sumr_230<= mulr_1_230 xor mulr_2_230;
sumr_231<= mulr_1_231 xor mulr_2_231;
sumr_232<= mulr_1_232 xor mulr_2_232;
sumr_233<= mulr_1_233 xor mulr_2_233;
sumr_234<= mulr_1_234 xor mulr_2_234;
sumr_235<= mulr_1_235 xor mulr_2_235;
sumr_236<= mulr_1_236 xor mulr_2_236;
sumr_237<= mulr_1_237 xor mulr_2_237;
sumr_238<= mulr_1_238 xor mulr_2_238;
sumr_239<= mulr_1_239 xor mulr_2_239;
sumr_240<= mulr_1_240 xor mulr_2_240;
sumr_241<= mulr_1_241 xor mulr_2_241;
sumr_242<= mulr_1_242 xor mulr_2_242;
sumr_243<= mulr_1_243 xor mulr_2_243;
sumr_244<= mulr_1_244 xor mulr_2_244;
sumr_245<= mulr_1_245 xor mulr_2_245;
sumr_246<= mulr_1_246 xor mulr_2_246;
sumr_247<= mulr_1_247 xor mulr_2_247;
sumr_248<= mulr_1_248 xor mulr_2_248;
sumr_249<= mulr_1_249 xor mulr_2_249;
sumr_250<= mulr_1_250 xor mulr_2_250;
sumr_251<= mulr_1_251 xor mulr_2_251;
sumr_252<= mulr_1_252 xor mulr_2_252;
sumr_253<= mulr_1_253 xor mulr_2_253;
sumr_254<= mulr_1_254 xor mulr_2_254;
sumr_255<= mulr_1_255 xor mulr_2_255;
sumr_256<= mulr_1_256 xor mulr_2_256;
sumr_257<= mulr_1_257 xor mulr_2_257;
sumr_258<= mulr_1_258 xor mulr_2_258;
sumr_259<= mulr_1_259 xor mulr_2_259;
sumr_260<= mulr_1_260 xor mulr_2_260;
sumr_261<= mulr_1_261 xor mulr_2_261;
sumr_262<= mulr_1_262 xor mulr_2_262;
sumr_263<= mulr_1_263 xor mulr_2_263;
sumr_264<= mulr_1_264 xor mulr_2_264;
sumr_265<= mulr_1_265 xor mulr_2_265;
sumr_266<= mulr_1_266 xor mulr_2_266;
sumr_267<= mulr_1_267 xor mulr_2_267;
sumr_268<= mulr_1_268 xor mulr_2_268;
sumr_269<= mulr_1_269 xor mulr_2_269;
sumr_270<= mulr_1_270 xor mulr_2_270;
sumr_271<= mulr_1_271 xor mulr_2_271;
sumr_272<= mulr_1_272 xor mulr_2_272;
sumr_273<= mulr_1_273 xor mulr_2_273;
sumr_274<= mulr_1_274 xor mulr_2_274;
sumr_275<= mulr_1_275 xor mulr_2_275;
sumr_276<= mulr_1_276 xor mulr_2_276;
sumr_277<= mulr_1_277 xor mulr_2_277;
sumr_278<= mulr_1_278 xor mulr_2_278;
sumr_279<= mulr_1_279 xor mulr_2_279;
sumr_280<= mulr_1_280 xor mulr_2_280;
sumr_281<= mulr_1_281 xor mulr_2_281;
sumr_282<= mulr_1_282 xor mulr_2_282;
sumr_283<= mulr_1_283 xor mulr_2_283;
sumr_284<= mulr_1_284 xor mulr_2_284;
sumr_285<= mulr_1_285 xor mulr_2_285;
sumr_286<= mulr_1_286 xor mulr_2_286;
sumr_287<= mulr_1_287 xor mulr_2_287;
sumr_288<= mulr_1_288 xor mulr_2_288;
sumr_289<= mulr_1_289 xor mulr_2_289;
sumr_290<= mulr_1_290 xor mulr_2_290;
sumr_291<= mulr_1_291 xor mulr_2_291;
sumr_292<= mulr_1_292 xor mulr_2_292;
sumr_293<= mulr_1_293 xor mulr_2_293;
sumr_294<= mulr_1_294 xor mulr_2_294;
sumr_295<= mulr_1_295 xor mulr_2_295;
sumr_296<= mulr_1_296 xor mulr_2_296;
sumr_297<= mulr_1_297 xor mulr_2_297;
sumr_298<= mulr_1_298 xor mulr_2_298;
sumr_299<= mulr_1_299 xor mulr_2_299;
sumr_300<= mulr_1_300 xor mulr_2_300;
sumr_301<= mulr_1_301 xor mulr_2_301;
sumr_302<= mulr_1_302 xor mulr_2_302;
sumr_303<= mulr_1_303 xor mulr_2_303;
sumr_304<= mulr_1_304 xor mulr_2_304;
sumr_305<= mulr_1_305 xor mulr_2_305;
sumr_306<= mulr_1_306 xor mulr_2_306;
sumr_307<= mulr_1_307 xor mulr_2_307;
sumr_308<= mulr_1_308 xor mulr_2_308;
sumr_309<= mulr_1_309 xor mulr_2_309;
sumr_310<= mulr_1_310 xor mulr_2_310;
sumr_311<= mulr_1_311 xor mulr_2_311;
sumr_312<= mulr_1_312 xor mulr_2_312;
sumr_313<= mulr_1_313 xor mulr_2_313;
sumr_314<= mulr_1_314 xor mulr_2_314;
sumr_315<= mulr_1_315 xor mulr_2_315;
sumr_316<= mulr_1_316 xor mulr_2_316;
sumr_317<= mulr_1_317 xor mulr_2_317;
sumr_318<= mulr_1_318 xor mulr_2_318;
sumr_319<= mulr_1_319 xor mulr_2_319;
sumr_320<= mulr_1_320 xor mulr_2_320;
sumr_321<= mulr_1_321 xor mulr_2_321;
sumr_322<= mulr_1_322 xor mulr_2_322;
sumr_323<= mulr_1_323 xor mulr_2_323;
sumr_324<= mulr_1_324 xor mulr_2_324;
sumr_325<= mulr_1_325 xor mulr_2_325;
sumr_326<= mulr_1_326 xor mulr_2_326;
sumr_327<= mulr_1_327 xor mulr_2_327;
sumr_328<= mulr_1_328 xor mulr_2_328;
sumr_329<= mulr_1_329 xor mulr_2_329;
sumr_330<= mulr_1_330 xor mulr_2_330;
sumr_331<= mulr_1_331 xor mulr_2_331;
sumr_332<= mulr_1_332 xor mulr_2_332;
sumr_333<= mulr_1_333 xor mulr_2_333;
sumr_334<= mulr_1_334 xor mulr_2_334;
sumr_335<= mulr_1_335 xor mulr_2_335;
sumr_336<= mulr_1_336 xor mulr_2_336;
sumr_337<= mulr_1_337 xor mulr_2_337;
sumr_338<= mulr_1_338 xor mulr_2_338;
sumr_339<= mulr_1_339 xor mulr_2_339;
sumr_340<= mulr_1_340 xor mulr_2_340;
sumr_341<= mulr_1_341 xor mulr_2_341;
sumr_342<= mulr_1_342 xor mulr_2_342;
sumr_343<= mulr_1_343 xor mulr_2_343;
sumr_344<= mulr_1_344 xor mulr_2_344;
sumr_345<= mulr_1_345 xor mulr_2_345;
sumr_346<= mulr_1_346 xor mulr_2_346;
sumr_347<= mulr_1_347 xor mulr_2_347;
sumr_348<= mulr_1_348 xor mulr_2_348;
sumr_349<= mulr_1_349 xor mulr_2_349;
sumr_350<= mulr_1_350 xor mulr_2_350;
sumr_351<= mulr_1_351 xor mulr_2_351;
sumr_352<= mulr_1_352 xor mulr_2_352;
sumr_353<= mulr_1_353 xor mulr_2_353;
sumr_354<= mulr_1_354 xor mulr_2_354;
sumr_355<= mulr_1_355 xor mulr_2_355;
sumr_356<= mulr_1_356 xor mulr_2_356;
sumr_357<= mulr_1_357 xor mulr_2_357;
sumr_358<= mulr_1_358 xor mulr_2_358;
sumr_359<= mulr_1_359 xor mulr_2_359;
sumr_360<= mulr_1_360 xor mulr_2_360;
sumr_361<= mulr_1_361 xor mulr_2_361;
sumr_362<= mulr_1_362 xor mulr_2_362;
sumr_363<= mulr_1_363 xor mulr_2_363;
sumr_364<= mulr_1_364 xor mulr_2_364;
sumr_365<= mulr_1_365 xor mulr_2_365;
sumr_366<= mulr_1_366 xor mulr_2_366;
sumr_367<= mulr_1_367 xor mulr_2_367;
sumr_368<= mulr_1_368 xor mulr_2_368;
sumr_369<= mulr_1_369 xor mulr_2_369;
sumr_370<= mulr_1_370 xor mulr_2_370;
sumr_371<= mulr_1_371 xor mulr_2_371;
sumr_372<= mulr_1_372 xor mulr_2_372;
sumr_373<= mulr_1_373 xor mulr_2_373;
sumr_374<= mulr_1_374 xor mulr_2_374;
sumr_375<= mulr_1_375 xor mulr_2_375;
sumr_376<= mulr_1_376 xor mulr_2_376;
sumr_377<= mulr_1_377 xor mulr_2_377;
sumr_378<= mulr_1_378 xor mulr_2_378;
sumr_379<= mulr_1_379 xor mulr_2_379;
sumr_380<= mulr_1_380 xor mulr_2_380;
sumr_381<= mulr_1_381 xor mulr_2_381;
sumr_382<= mulr_1_382 xor mulr_2_382;
sumr_383<= mulr_1_383 xor mulr_2_383;
sumr_384<= mulr_1_384 xor mulr_2_384;
sumr_385<= mulr_1_385 xor mulr_2_385;
sumr_386<= mulr_1_386 xor mulr_2_386;
sumr_387<= mulr_1_387 xor mulr_2_387;
sumr_388<= mulr_1_388 xor mulr_2_388;
sumr_389<= mulr_1_389 xor mulr_2_389;
sumr_390<= mulr_1_390 xor mulr_2_390;
sumr_391<= mulr_1_391 xor mulr_2_391;
sumr_392<= mulr_1_392 xor mulr_2_392;
sumr_393<= mulr_1_393 xor mulr_2_393;
sumr_394<= mulr_1_394 xor mulr_2_394;
sumr_395<= mulr_1_395 xor mulr_2_395;
sumr_396<= mulr_1_396 xor mulr_2_396;
sumr_397<= mulr_1_397 xor mulr_2_397;
sumr_398<= mulr_1_398 xor mulr_2_398;
sumr_399<= mulr_1_399 xor mulr_2_399;
sumr_400<= mulr_1_400 xor mulr_2_400;
sumr_401<= mulr_1_401 xor mulr_2_401;
sumr_402<= mulr_1_402 xor mulr_2_402;
sumr_403<= mulr_1_403 xor mulr_2_403;
sumr_404<= mulr_1_404 xor mulr_2_404;
sumr_405<= mulr_1_405 xor mulr_2_405;
sumr_406<= mulr_1_406 xor mulr_2_406;
sumr_407<= mulr_1_407 xor mulr_2_407;
sumr_408<= mulr_1_408 xor mulr_2_408;
sumr_409<= mulr_1_409 xor mulr_2_409;
sumr_410<= mulr_1_410 xor mulr_2_410;
sumr_411<= mulr_1_411 xor mulr_2_411;
sumr_412<= mulr_1_412 xor mulr_2_412;
sumr_413<= mulr_1_413 xor mulr_2_413;
sumr_414<= mulr_1_414 xor mulr_2_414;
sumr_415<= mulr_1_415 xor mulr_2_415;
sumr_416<= mulr_1_416 xor mulr_2_416;
sumr_417<= mulr_1_417 xor mulr_2_417;
sumr_418<= mulr_1_418 xor mulr_2_418;
sumr_419<= mulr_1_419 xor mulr_2_419;
sumr_420<= mulr_1_420 xor mulr_2_420;
sumr_421<= mulr_1_421 xor mulr_2_421;
sumr_422<= mulr_1_422 xor mulr_2_422;
sumr_423<= mulr_1_423 xor mulr_2_423;
sumr_424<= mulr_1_424 xor mulr_2_424;
sumr_425<= mulr_1_425 xor mulr_2_425;
sumr_426<= mulr_1_426 xor mulr_2_426;
sumr_427<= mulr_1_427 xor mulr_2_427;
sumr_428<= mulr_1_428 xor mulr_2_428;
sumr_429<= mulr_1_429 xor mulr_2_429;
sumr_430<= mulr_1_430 xor mulr_2_430;
sumr_431<= mulr_1_431 xor mulr_2_431;
sumr_432<= mulr_1_432 xor mulr_2_432;
sumr_433<= mulr_1_433 xor mulr_2_433;
sumr_434<= mulr_1_434 xor mulr_2_434;
sumr_435<= mulr_1_435 xor mulr_2_435;
sumr_436<= mulr_1_436 xor mulr_2_436;
sumr_437<= mulr_1_437 xor mulr_2_437;
sumr_438<= mulr_1_438 xor mulr_2_438;
sumr_439<= mulr_1_439 xor mulr_2_439;
sumr_440<= mulr_1_440 xor mulr_2_440;
sumr_441<= mulr_1_441 xor mulr_2_441;
sumr_442<= mulr_1_442 xor mulr_2_442;
sumr_443<= mulr_1_443 xor mulr_2_443;
sumr_444<= mulr_1_444 xor mulr_2_444;
sumr_445<= mulr_1_445 xor mulr_2_445;
sumr_446<= mulr_1_446 xor mulr_2_446;
sumr_447<= mulr_1_447 xor mulr_2_447;
sumr_448<= mulr_1_448 xor mulr_2_448;
sumr_449<= mulr_1_449 xor mulr_2_449;
sumr_450<= mulr_1_450 xor mulr_2_450;
sumr_451<= mulr_1_451 xor mulr_2_451;
sumr_452<= mulr_1_452 xor mulr_2_452;
sumr_453<= mulr_1_453 xor mulr_2_453;
sumr_454<= mulr_1_454 xor mulr_2_454;
sumr_455<= mulr_1_455 xor mulr_2_455;
sumr_456<= mulr_1_456 xor mulr_2_456;
sumr_457<= mulr_1_457 xor mulr_2_457;
sumr_458<= mulr_1_458 xor mulr_2_458;
sumr_459<= mulr_1_459 xor mulr_2_459;
sumr_460<= mulr_1_460 xor mulr_2_460;
sumr_461<= mulr_1_461 xor mulr_2_461;
sumr_462<= mulr_1_462 xor mulr_2_462;
sumr_463<= mulr_1_463 xor mulr_2_463;
sumr_464<= mulr_1_464 xor mulr_2_464;
sumr_465<= mulr_1_465 xor mulr_2_465;
sumr_466<= mulr_1_466 xor mulr_2_466;
sumr_467<= mulr_1_467 xor mulr_2_467;
sumr_468<= mulr_1_468 xor mulr_2_468;
sumr_469<= mulr_1_469 xor mulr_2_469;
sumr_470<= mulr_1_470 xor mulr_2_470;
sumr_471<= mulr_1_471 xor mulr_2_471;
sumr_472<= mulr_1_472 xor mulr_2_472;
sumr_473<= mulr_1_473 xor mulr_2_473;
sumr_474<= mulr_1_474 xor mulr_2_474;
sumr_475<= mulr_1_475 xor mulr_2_475;
sumr_476<= mulr_1_476 xor mulr_2_476;
sumr_477<= mulr_1_477 xor mulr_2_477;
sumr_478<= mulr_1_478 xor mulr_2_478;
sumr_479<= mulr_1_479 xor mulr_2_479;
sumr_480<= mulr_1_480 xor mulr_2_480;
sumr_481<= mulr_1_481 xor mulr_2_481;
sumr_482<= mulr_1_482 xor mulr_2_482;
sumr_483<= mulr_1_483 xor mulr_2_483;
sumr_484<= mulr_1_484 xor mulr_2_484;
sumr_485<= mulr_1_485 xor mulr_2_485;
sumr_486<= mulr_1_486 xor mulr_2_486;
sumr_487<= mulr_1_487 xor mulr_2_487;
sumr_488<= mulr_1_488 xor mulr_2_488;
sumr_489<= mulr_1_489 xor mulr_2_489;
sumr_490<= mulr_1_490 xor mulr_2_490;
sumr_491<= mulr_1_491 xor mulr_2_491;
sumr_492<= mulr_1_492 xor mulr_2_492;
sumr_493<= mulr_1_493 xor mulr_2_493;
sumr_494<= mulr_1_494 xor mulr_2_494;
sumr_495<= mulr_1_495 xor mulr_2_495;
sumr_496<= mulr_1_496 xor mulr_2_496;
sumr_497<= mulr_1_497 xor mulr_2_497;
sumr_498<= mulr_1_498 xor mulr_2_498;
sumr_499<= mulr_1_499 xor mulr_2_499;
sumr_500<= mulr_1_500 xor mulr_2_500;
sumr_501<= mulr_1_501 xor mulr_2_501;
sumr_502<= mulr_1_502 xor mulr_2_502;
sumr_503<= mulr_1_503 xor mulr_2_503;
sumr_504<= mulr_1_504 xor mulr_2_504;
sumr_505<= mulr_1_505 xor mulr_2_505;
sumr_506<= mulr_1_506 xor mulr_2_506;
sumr_507<= mulr_1_507 xor mulr_2_507;
sumr_508<= mulr_1_508 xor mulr_2_508;
sumr_509<= mulr_1_509 xor mulr_2_509;
sumr_510<= mulr_1_510 xor mulr_2_510;
sumr_511<= mulr_1_511 xor mulr_2_511;
E(510)<=not ( sumr_1(0) or sumr_1(1) or sumr_1(2) or sumr_1(3) or sumr_1(4) or sumr_1(5) or sumr_1(6) or sumr_1(7) or sumr_1(8));
E(509)<=not ( sumr_2(0) or sumr_2(1) or sumr_2(2) or sumr_2(3) or sumr_2(4) or sumr_2(5) or sumr_2(6) or sumr_2(7) or sumr_2(8));
E(508)<=not ( sumr_3(0) or sumr_3(1) or sumr_3(2) or sumr_3(3) or sumr_3(4) or sumr_3(5) or sumr_3(6) or sumr_3(7) or sumr_3(8));
E(507)<=not ( sumr_4(0) or sumr_4(1) or sumr_4(2) or sumr_4(3) or sumr_4(4) or sumr_4(5) or sumr_4(6) or sumr_4(7) or sumr_4(8));
E(506)<=not ( sumr_5(0) or sumr_5(1) or sumr_5(2) or sumr_5(3) or sumr_5(4) or sumr_5(5) or sumr_5(6) or sumr_5(7) or sumr_5(8));
E(505)<=not ( sumr_6(0) or sumr_6(1) or sumr_6(2) or sumr_6(3) or sumr_6(4) or sumr_6(5) or sumr_6(6) or sumr_6(7) or sumr_6(8));
E(504)<=not ( sumr_7(0) or sumr_7(1) or sumr_7(2) or sumr_7(3) or sumr_7(4) or sumr_7(5) or sumr_7(6) or sumr_7(7) or sumr_7(8));
E(503)<=not ( sumr_8(0) or sumr_8(1) or sumr_8(2) or sumr_8(3) or sumr_8(4) or sumr_8(5) or sumr_8(6) or sumr_8(7) or sumr_8(8));
E(502)<=not ( sumr_9(0) or sumr_9(1) or sumr_9(2) or sumr_9(3) or sumr_9(4) or sumr_9(5) or sumr_9(6) or sumr_9(7) or sumr_9(8));
E(501)<=not ( sumr_10(0) or sumr_10(1) or sumr_10(2) or sumr_10(3) or sumr_10(4) or sumr_10(5) or sumr_10(6) or sumr_10(7) or sumr_10(8));
E(500)<=not ( sumr_11(0) or sumr_11(1) or sumr_11(2) or sumr_11(3) or sumr_11(4) or sumr_11(5) or sumr_11(6) or sumr_11(7) or sumr_11(8));
E(499)<=not ( sumr_12(0) or sumr_12(1) or sumr_12(2) or sumr_12(3) or sumr_12(4) or sumr_12(5) or sumr_12(6) or sumr_12(7) or sumr_12(8));
E(498)<=not ( sumr_13(0) or sumr_13(1) or sumr_13(2) or sumr_13(3) or sumr_13(4) or sumr_13(5) or sumr_13(6) or sumr_13(7) or sumr_13(8));
E(497)<=not ( sumr_14(0) or sumr_14(1) or sumr_14(2) or sumr_14(3) or sumr_14(4) or sumr_14(5) or sumr_14(6) or sumr_14(7) or sumr_14(8));
E(496)<=not ( sumr_15(0) or sumr_15(1) or sumr_15(2) or sumr_15(3) or sumr_15(4) or sumr_15(5) or sumr_15(6) or sumr_15(7) or sumr_15(8));
E(495)<=not ( sumr_16(0) or sumr_16(1) or sumr_16(2) or sumr_16(3) or sumr_16(4) or sumr_16(5) or sumr_16(6) or sumr_16(7) or sumr_16(8));
E(494)<=not ( sumr_17(0) or sumr_17(1) or sumr_17(2) or sumr_17(3) or sumr_17(4) or sumr_17(5) or sumr_17(6) or sumr_17(7) or sumr_17(8));
E(493)<=not ( sumr_18(0) or sumr_18(1) or sumr_18(2) or sumr_18(3) or sumr_18(4) or sumr_18(5) or sumr_18(6) or sumr_18(7) or sumr_18(8));
E(492)<=not ( sumr_19(0) or sumr_19(1) or sumr_19(2) or sumr_19(3) or sumr_19(4) or sumr_19(5) or sumr_19(6) or sumr_19(7) or sumr_19(8));
E(491)<=not ( sumr_20(0) or sumr_20(1) or sumr_20(2) or sumr_20(3) or sumr_20(4) or sumr_20(5) or sumr_20(6) or sumr_20(7) or sumr_20(8));
E(490)<=not ( sumr_21(0) or sumr_21(1) or sumr_21(2) or sumr_21(3) or sumr_21(4) or sumr_21(5) or sumr_21(6) or sumr_21(7) or sumr_21(8));
E(489)<=not ( sumr_22(0) or sumr_22(1) or sumr_22(2) or sumr_22(3) or sumr_22(4) or sumr_22(5) or sumr_22(6) or sumr_22(7) or sumr_22(8));
E(488)<=not ( sumr_23(0) or sumr_23(1) or sumr_23(2) or sumr_23(3) or sumr_23(4) or sumr_23(5) or sumr_23(6) or sumr_23(7) or sumr_23(8));
E(487)<=not ( sumr_24(0) or sumr_24(1) or sumr_24(2) or sumr_24(3) or sumr_24(4) or sumr_24(5) or sumr_24(6) or sumr_24(7) or sumr_24(8));
E(486)<=not ( sumr_25(0) or sumr_25(1) or sumr_25(2) or sumr_25(3) or sumr_25(4) or sumr_25(5) or sumr_25(6) or sumr_25(7) or sumr_25(8));
E(485)<=not ( sumr_26(0) or sumr_26(1) or sumr_26(2) or sumr_26(3) or sumr_26(4) or sumr_26(5) or sumr_26(6) or sumr_26(7) or sumr_26(8));
E(484)<=not ( sumr_27(0) or sumr_27(1) or sumr_27(2) or sumr_27(3) or sumr_27(4) or sumr_27(5) or sumr_27(6) or sumr_27(7) or sumr_27(8));
E(483)<=not ( sumr_28(0) or sumr_28(1) or sumr_28(2) or sumr_28(3) or sumr_28(4) or sumr_28(5) or sumr_28(6) or sumr_28(7) or sumr_28(8));
E(482)<=not ( sumr_29(0) or sumr_29(1) or sumr_29(2) or sumr_29(3) or sumr_29(4) or sumr_29(5) or sumr_29(6) or sumr_29(7) or sumr_29(8));
E(481)<=not ( sumr_30(0) or sumr_30(1) or sumr_30(2) or sumr_30(3) or sumr_30(4) or sumr_30(5) or sumr_30(6) or sumr_30(7) or sumr_30(8));
E(480)<=not ( sumr_31(0) or sumr_31(1) or sumr_31(2) or sumr_31(3) or sumr_31(4) or sumr_31(5) or sumr_31(6) or sumr_31(7) or sumr_31(8));
E(479)<=not ( sumr_32(0) or sumr_32(1) or sumr_32(2) or sumr_32(3) or sumr_32(4) or sumr_32(5) or sumr_32(6) or sumr_32(7) or sumr_32(8));
E(478)<=not ( sumr_33(0) or sumr_33(1) or sumr_33(2) or sumr_33(3) or sumr_33(4) or sumr_33(5) or sumr_33(6) or sumr_33(7) or sumr_33(8));
E(477)<=not ( sumr_34(0) or sumr_34(1) or sumr_34(2) or sumr_34(3) or sumr_34(4) or sumr_34(5) or sumr_34(6) or sumr_34(7) or sumr_34(8));
E(476)<=not ( sumr_35(0) or sumr_35(1) or sumr_35(2) or sumr_35(3) or sumr_35(4) or sumr_35(5) or sumr_35(6) or sumr_35(7) or sumr_35(8));
E(475)<=not ( sumr_36(0) or sumr_36(1) or sumr_36(2) or sumr_36(3) or sumr_36(4) or sumr_36(5) or sumr_36(6) or sumr_36(7) or sumr_36(8));
E(474)<=not ( sumr_37(0) or sumr_37(1) or sumr_37(2) or sumr_37(3) or sumr_37(4) or sumr_37(5) or sumr_37(6) or sumr_37(7) or sumr_37(8));
E(473)<=not ( sumr_38(0) or sumr_38(1) or sumr_38(2) or sumr_38(3) or sumr_38(4) or sumr_38(5) or sumr_38(6) or sumr_38(7) or sumr_38(8));
E(472)<=not ( sumr_39(0) or sumr_39(1) or sumr_39(2) or sumr_39(3) or sumr_39(4) or sumr_39(5) or sumr_39(6) or sumr_39(7) or sumr_39(8));
E(471)<=not ( sumr_40(0) or sumr_40(1) or sumr_40(2) or sumr_40(3) or sumr_40(4) or sumr_40(5) or sumr_40(6) or sumr_40(7) or sumr_40(8));
E(470)<=not ( sumr_41(0) or sumr_41(1) or sumr_41(2) or sumr_41(3) or sumr_41(4) or sumr_41(5) or sumr_41(6) or sumr_41(7) or sumr_41(8));
E(469)<=not ( sumr_42(0) or sumr_42(1) or sumr_42(2) or sumr_42(3) or sumr_42(4) or sumr_42(5) or sumr_42(6) or sumr_42(7) or sumr_42(8));
E(468)<=not ( sumr_43(0) or sumr_43(1) or sumr_43(2) or sumr_43(3) or sumr_43(4) or sumr_43(5) or sumr_43(6) or sumr_43(7) or sumr_43(8));
E(467)<=not ( sumr_44(0) or sumr_44(1) or sumr_44(2) or sumr_44(3) or sumr_44(4) or sumr_44(5) or sumr_44(6) or sumr_44(7) or sumr_44(8));
E(466)<=not ( sumr_45(0) or sumr_45(1) or sumr_45(2) or sumr_45(3) or sumr_45(4) or sumr_45(5) or sumr_45(6) or sumr_45(7) or sumr_45(8));
E(465)<=not ( sumr_46(0) or sumr_46(1) or sumr_46(2) or sumr_46(3) or sumr_46(4) or sumr_46(5) or sumr_46(6) or sumr_46(7) or sumr_46(8));
E(464)<=not ( sumr_47(0) or sumr_47(1) or sumr_47(2) or sumr_47(3) or sumr_47(4) or sumr_47(5) or sumr_47(6) or sumr_47(7) or sumr_47(8));
E(463)<=not ( sumr_48(0) or sumr_48(1) or sumr_48(2) or sumr_48(3) or sumr_48(4) or sumr_48(5) or sumr_48(6) or sumr_48(7) or sumr_48(8));
E(462)<=not ( sumr_49(0) or sumr_49(1) or sumr_49(2) or sumr_49(3) or sumr_49(4) or sumr_49(5) or sumr_49(6) or sumr_49(7) or sumr_49(8));
E(461)<=not ( sumr_50(0) or sumr_50(1) or sumr_50(2) or sumr_50(3) or sumr_50(4) or sumr_50(5) or sumr_50(6) or sumr_50(7) or sumr_50(8));
E(460)<=not ( sumr_51(0) or sumr_51(1) or sumr_51(2) or sumr_51(3) or sumr_51(4) or sumr_51(5) or sumr_51(6) or sumr_51(7) or sumr_51(8));
E(459)<=not ( sumr_52(0) or sumr_52(1) or sumr_52(2) or sumr_52(3) or sumr_52(4) or sumr_52(5) or sumr_52(6) or sumr_52(7) or sumr_52(8));
E(458)<=not ( sumr_53(0) or sumr_53(1) or sumr_53(2) or sumr_53(3) or sumr_53(4) or sumr_53(5) or sumr_53(6) or sumr_53(7) or sumr_53(8));
E(457)<=not ( sumr_54(0) or sumr_54(1) or sumr_54(2) or sumr_54(3) or sumr_54(4) or sumr_54(5) or sumr_54(6) or sumr_54(7) or sumr_54(8));
E(456)<=not ( sumr_55(0) or sumr_55(1) or sumr_55(2) or sumr_55(3) or sumr_55(4) or sumr_55(5) or sumr_55(6) or sumr_55(7) or sumr_55(8));
E(455)<=not ( sumr_56(0) or sumr_56(1) or sumr_56(2) or sumr_56(3) or sumr_56(4) or sumr_56(5) or sumr_56(6) or sumr_56(7) or sumr_56(8));
E(454)<=not ( sumr_57(0) or sumr_57(1) or sumr_57(2) or sumr_57(3) or sumr_57(4) or sumr_57(5) or sumr_57(6) or sumr_57(7) or sumr_57(8));
E(453)<=not ( sumr_58(0) or sumr_58(1) or sumr_58(2) or sumr_58(3) or sumr_58(4) or sumr_58(5) or sumr_58(6) or sumr_58(7) or sumr_58(8));
E(452)<=not ( sumr_59(0) or sumr_59(1) or sumr_59(2) or sumr_59(3) or sumr_59(4) or sumr_59(5) or sumr_59(6) or sumr_59(7) or sumr_59(8));
E(451)<=not ( sumr_60(0) or sumr_60(1) or sumr_60(2) or sumr_60(3) or sumr_60(4) or sumr_60(5) or sumr_60(6) or sumr_60(7) or sumr_60(8));
E(450)<=not ( sumr_61(0) or sumr_61(1) or sumr_61(2) or sumr_61(3) or sumr_61(4) or sumr_61(5) or sumr_61(6) or sumr_61(7) or sumr_61(8));
E(449)<=not ( sumr_62(0) or sumr_62(1) or sumr_62(2) or sumr_62(3) or sumr_62(4) or sumr_62(5) or sumr_62(6) or sumr_62(7) or sumr_62(8));
E(448)<=not ( sumr_63(0) or sumr_63(1) or sumr_63(2) or sumr_63(3) or sumr_63(4) or sumr_63(5) or sumr_63(6) or sumr_63(7) or sumr_63(8));
E(447)<=not ( sumr_64(0) or sumr_64(1) or sumr_64(2) or sumr_64(3) or sumr_64(4) or sumr_64(5) or sumr_64(6) or sumr_64(7) or sumr_64(8));
E(446)<=not ( sumr_65(0) or sumr_65(1) or sumr_65(2) or sumr_65(3) or sumr_65(4) or sumr_65(5) or sumr_65(6) or sumr_65(7) or sumr_65(8));
E(445)<=not ( sumr_66(0) or sumr_66(1) or sumr_66(2) or sumr_66(3) or sumr_66(4) or sumr_66(5) or sumr_66(6) or sumr_66(7) or sumr_66(8));
E(444)<=not ( sumr_67(0) or sumr_67(1) or sumr_67(2) or sumr_67(3) or sumr_67(4) or sumr_67(5) or sumr_67(6) or sumr_67(7) or sumr_67(8));
E(443)<=not ( sumr_68(0) or sumr_68(1) or sumr_68(2) or sumr_68(3) or sumr_68(4) or sumr_68(5) or sumr_68(6) or sumr_68(7) or sumr_68(8));
E(442)<=not ( sumr_69(0) or sumr_69(1) or sumr_69(2) or sumr_69(3) or sumr_69(4) or sumr_69(5) or sumr_69(6) or sumr_69(7) or sumr_69(8));
E(441)<=not ( sumr_70(0) or sumr_70(1) or sumr_70(2) or sumr_70(3) or sumr_70(4) or sumr_70(5) or sumr_70(6) or sumr_70(7) or sumr_70(8));
E(440)<=not ( sumr_71(0) or sumr_71(1) or sumr_71(2) or sumr_71(3) or sumr_71(4) or sumr_71(5) or sumr_71(6) or sumr_71(7) or sumr_71(8));
E(439)<=not ( sumr_72(0) or sumr_72(1) or sumr_72(2) or sumr_72(3) or sumr_72(4) or sumr_72(5) or sumr_72(6) or sumr_72(7) or sumr_72(8));
E(438)<=not ( sumr_73(0) or sumr_73(1) or sumr_73(2) or sumr_73(3) or sumr_73(4) or sumr_73(5) or sumr_73(6) or sumr_73(7) or sumr_73(8));
E(437)<=not ( sumr_74(0) or sumr_74(1) or sumr_74(2) or sumr_74(3) or sumr_74(4) or sumr_74(5) or sumr_74(6) or sumr_74(7) or sumr_74(8));
E(436)<=not ( sumr_75(0) or sumr_75(1) or sumr_75(2) or sumr_75(3) or sumr_75(4) or sumr_75(5) or sumr_75(6) or sumr_75(7) or sumr_75(8));
E(435)<=not ( sumr_76(0) or sumr_76(1) or sumr_76(2) or sumr_76(3) or sumr_76(4) or sumr_76(5) or sumr_76(6) or sumr_76(7) or sumr_76(8));
E(434)<=not ( sumr_77(0) or sumr_77(1) or sumr_77(2) or sumr_77(3) or sumr_77(4) or sumr_77(5) or sumr_77(6) or sumr_77(7) or sumr_77(8));
E(433)<=not ( sumr_78(0) or sumr_78(1) or sumr_78(2) or sumr_78(3) or sumr_78(4) or sumr_78(5) or sumr_78(6) or sumr_78(7) or sumr_78(8));
E(432)<=not ( sumr_79(0) or sumr_79(1) or sumr_79(2) or sumr_79(3) or sumr_79(4) or sumr_79(5) or sumr_79(6) or sumr_79(7) or sumr_79(8));
E(431)<=not ( sumr_80(0) or sumr_80(1) or sumr_80(2) or sumr_80(3) or sumr_80(4) or sumr_80(5) or sumr_80(6) or sumr_80(7) or sumr_80(8));
E(430)<=not ( sumr_81(0) or sumr_81(1) or sumr_81(2) or sumr_81(3) or sumr_81(4) or sumr_81(5) or sumr_81(6) or sumr_81(7) or sumr_81(8));
E(429)<=not ( sumr_82(0) or sumr_82(1) or sumr_82(2) or sumr_82(3) or sumr_82(4) or sumr_82(5) or sumr_82(6) or sumr_82(7) or sumr_82(8));
E(428)<=not ( sumr_83(0) or sumr_83(1) or sumr_83(2) or sumr_83(3) or sumr_83(4) or sumr_83(5) or sumr_83(6) or sumr_83(7) or sumr_83(8));
E(427)<=not ( sumr_84(0) or sumr_84(1) or sumr_84(2) or sumr_84(3) or sumr_84(4) or sumr_84(5) or sumr_84(6) or sumr_84(7) or sumr_84(8));
E(426)<=not ( sumr_85(0) or sumr_85(1) or sumr_85(2) or sumr_85(3) or sumr_85(4) or sumr_85(5) or sumr_85(6) or sumr_85(7) or sumr_85(8));
E(425)<=not ( sumr_86(0) or sumr_86(1) or sumr_86(2) or sumr_86(3) or sumr_86(4) or sumr_86(5) or sumr_86(6) or sumr_86(7) or sumr_86(8));
E(424)<=not ( sumr_87(0) or sumr_87(1) or sumr_87(2) or sumr_87(3) or sumr_87(4) or sumr_87(5) or sumr_87(6) or sumr_87(7) or sumr_87(8));
E(423)<=not ( sumr_88(0) or sumr_88(1) or sumr_88(2) or sumr_88(3) or sumr_88(4) or sumr_88(5) or sumr_88(6) or sumr_88(7) or sumr_88(8));
E(422)<=not ( sumr_89(0) or sumr_89(1) or sumr_89(2) or sumr_89(3) or sumr_89(4) or sumr_89(5) or sumr_89(6) or sumr_89(7) or sumr_89(8));
E(421)<=not ( sumr_90(0) or sumr_90(1) or sumr_90(2) or sumr_90(3) or sumr_90(4) or sumr_90(5) or sumr_90(6) or sumr_90(7) or sumr_90(8));
E(420)<=not ( sumr_91(0) or sumr_91(1) or sumr_91(2) or sumr_91(3) or sumr_91(4) or sumr_91(5) or sumr_91(6) or sumr_91(7) or sumr_91(8));
E(419)<=not ( sumr_92(0) or sumr_92(1) or sumr_92(2) or sumr_92(3) or sumr_92(4) or sumr_92(5) or sumr_92(6) or sumr_92(7) or sumr_92(8));
E(418)<=not ( sumr_93(0) or sumr_93(1) or sumr_93(2) or sumr_93(3) or sumr_93(4) or sumr_93(5) or sumr_93(6) or sumr_93(7) or sumr_93(8));
E(417)<=not ( sumr_94(0) or sumr_94(1) or sumr_94(2) or sumr_94(3) or sumr_94(4) or sumr_94(5) or sumr_94(6) or sumr_94(7) or sumr_94(8));
E(416)<=not ( sumr_95(0) or sumr_95(1) or sumr_95(2) or sumr_95(3) or sumr_95(4) or sumr_95(5) or sumr_95(6) or sumr_95(7) or sumr_95(8));
E(415)<=not ( sumr_96(0) or sumr_96(1) or sumr_96(2) or sumr_96(3) or sumr_96(4) or sumr_96(5) or sumr_96(6) or sumr_96(7) or sumr_96(8));
E(414)<=not ( sumr_97(0) or sumr_97(1) or sumr_97(2) or sumr_97(3) or sumr_97(4) or sumr_97(5) or sumr_97(6) or sumr_97(7) or sumr_97(8));
E(413)<=not ( sumr_98(0) or sumr_98(1) or sumr_98(2) or sumr_98(3) or sumr_98(4) or sumr_98(5) or sumr_98(6) or sumr_98(7) or sumr_98(8));
E(412)<=not ( sumr_99(0) or sumr_99(1) or sumr_99(2) or sumr_99(3) or sumr_99(4) or sumr_99(5) or sumr_99(6) or sumr_99(7) or sumr_99(8));
E(411)<=not ( sumr_100(0) or sumr_100(1) or sumr_100(2) or sumr_100(3) or sumr_100(4) or sumr_100(5) or sumr_100(6) or sumr_100(7) or sumr_100(8));
E(410)<=not ( sumr_101(0) or sumr_101(1) or sumr_101(2) or sumr_101(3) or sumr_101(4) or sumr_101(5) or sumr_101(6) or sumr_101(7) or sumr_101(8));
E(409)<=not ( sumr_102(0) or sumr_102(1) or sumr_102(2) or sumr_102(3) or sumr_102(4) or sumr_102(5) or sumr_102(6) or sumr_102(7) or sumr_102(8));
E(408)<=not ( sumr_103(0) or sumr_103(1) or sumr_103(2) or sumr_103(3) or sumr_103(4) or sumr_103(5) or sumr_103(6) or sumr_103(7) or sumr_103(8));
E(407)<=not ( sumr_104(0) or sumr_104(1) or sumr_104(2) or sumr_104(3) or sumr_104(4) or sumr_104(5) or sumr_104(6) or sumr_104(7) or sumr_104(8));
E(406)<=not ( sumr_105(0) or sumr_105(1) or sumr_105(2) or sumr_105(3) or sumr_105(4) or sumr_105(5) or sumr_105(6) or sumr_105(7) or sumr_105(8));
E(405)<=not ( sumr_106(0) or sumr_106(1) or sumr_106(2) or sumr_106(3) or sumr_106(4) or sumr_106(5) or sumr_106(6) or sumr_106(7) or sumr_106(8));
E(404)<=not ( sumr_107(0) or sumr_107(1) or sumr_107(2) or sumr_107(3) or sumr_107(4) or sumr_107(5) or sumr_107(6) or sumr_107(7) or sumr_107(8));
E(403)<=not ( sumr_108(0) or sumr_108(1) or sumr_108(2) or sumr_108(3) or sumr_108(4) or sumr_108(5) or sumr_108(6) or sumr_108(7) or sumr_108(8));
E(402)<=not ( sumr_109(0) or sumr_109(1) or sumr_109(2) or sumr_109(3) or sumr_109(4) or sumr_109(5) or sumr_109(6) or sumr_109(7) or sumr_109(8));
E(401)<=not ( sumr_110(0) or sumr_110(1) or sumr_110(2) or sumr_110(3) or sumr_110(4) or sumr_110(5) or sumr_110(6) or sumr_110(7) or sumr_110(8));
E(400)<=not ( sumr_111(0) or sumr_111(1) or sumr_111(2) or sumr_111(3) or sumr_111(4) or sumr_111(5) or sumr_111(6) or sumr_111(7) or sumr_111(8));
E(399)<=not ( sumr_112(0) or sumr_112(1) or sumr_112(2) or sumr_112(3) or sumr_112(4) or sumr_112(5) or sumr_112(6) or sumr_112(7) or sumr_112(8));
E(398)<=not ( sumr_113(0) or sumr_113(1) or sumr_113(2) or sumr_113(3) or sumr_113(4) or sumr_113(5) or sumr_113(6) or sumr_113(7) or sumr_113(8));
E(397)<=not ( sumr_114(0) or sumr_114(1) or sumr_114(2) or sumr_114(3) or sumr_114(4) or sumr_114(5) or sumr_114(6) or sumr_114(7) or sumr_114(8));
E(396)<=not ( sumr_115(0) or sumr_115(1) or sumr_115(2) or sumr_115(3) or sumr_115(4) or sumr_115(5) or sumr_115(6) or sumr_115(7) or sumr_115(8));
E(395)<=not ( sumr_116(0) or sumr_116(1) or sumr_116(2) or sumr_116(3) or sumr_116(4) or sumr_116(5) or sumr_116(6) or sumr_116(7) or sumr_116(8));
E(394)<=not ( sumr_117(0) or sumr_117(1) or sumr_117(2) or sumr_117(3) or sumr_117(4) or sumr_117(5) or sumr_117(6) or sumr_117(7) or sumr_117(8));
E(393)<=not ( sumr_118(0) or sumr_118(1) or sumr_118(2) or sumr_118(3) or sumr_118(4) or sumr_118(5) or sumr_118(6) or sumr_118(7) or sumr_118(8));
E(392)<=not ( sumr_119(0) or sumr_119(1) or sumr_119(2) or sumr_119(3) or sumr_119(4) or sumr_119(5) or sumr_119(6) or sumr_119(7) or sumr_119(8));
E(391)<=not ( sumr_120(0) or sumr_120(1) or sumr_120(2) or sumr_120(3) or sumr_120(4) or sumr_120(5) or sumr_120(6) or sumr_120(7) or sumr_120(8));
E(390)<=not ( sumr_121(0) or sumr_121(1) or sumr_121(2) or sumr_121(3) or sumr_121(4) or sumr_121(5) or sumr_121(6) or sumr_121(7) or sumr_121(8));
E(389)<=not ( sumr_122(0) or sumr_122(1) or sumr_122(2) or sumr_122(3) or sumr_122(4) or sumr_122(5) or sumr_122(6) or sumr_122(7) or sumr_122(8));
E(388)<=not ( sumr_123(0) or sumr_123(1) or sumr_123(2) or sumr_123(3) or sumr_123(4) or sumr_123(5) or sumr_123(6) or sumr_123(7) or sumr_123(8));
E(387)<=not ( sumr_124(0) or sumr_124(1) or sumr_124(2) or sumr_124(3) or sumr_124(4) or sumr_124(5) or sumr_124(6) or sumr_124(7) or sumr_124(8));
E(386)<=not ( sumr_125(0) or sumr_125(1) or sumr_125(2) or sumr_125(3) or sumr_125(4) or sumr_125(5) or sumr_125(6) or sumr_125(7) or sumr_125(8));
E(385)<=not ( sumr_126(0) or sumr_126(1) or sumr_126(2) or sumr_126(3) or sumr_126(4) or sumr_126(5) or sumr_126(6) or sumr_126(7) or sumr_126(8));
E(384)<=not ( sumr_127(0) or sumr_127(1) or sumr_127(2) or sumr_127(3) or sumr_127(4) or sumr_127(5) or sumr_127(6) or sumr_127(7) or sumr_127(8));
E(383)<=not ( sumr_128(0) or sumr_128(1) or sumr_128(2) or sumr_128(3) or sumr_128(4) or sumr_128(5) or sumr_128(6) or sumr_128(7) or sumr_128(8));
E(382)<=not ( sumr_129(0) or sumr_129(1) or sumr_129(2) or sumr_129(3) or sumr_129(4) or sumr_129(5) or sumr_129(6) or sumr_129(7) or sumr_129(8));
E(381)<=not ( sumr_130(0) or sumr_130(1) or sumr_130(2) or sumr_130(3) or sumr_130(4) or sumr_130(5) or sumr_130(6) or sumr_130(7) or sumr_130(8));
E(380)<=not ( sumr_131(0) or sumr_131(1) or sumr_131(2) or sumr_131(3) or sumr_131(4) or sumr_131(5) or sumr_131(6) or sumr_131(7) or sumr_131(8));
E(379)<=not ( sumr_132(0) or sumr_132(1) or sumr_132(2) or sumr_132(3) or sumr_132(4) or sumr_132(5) or sumr_132(6) or sumr_132(7) or sumr_132(8));
E(378)<=not ( sumr_133(0) or sumr_133(1) or sumr_133(2) or sumr_133(3) or sumr_133(4) or sumr_133(5) or sumr_133(6) or sumr_133(7) or sumr_133(8));
E(377)<=not ( sumr_134(0) or sumr_134(1) or sumr_134(2) or sumr_134(3) or sumr_134(4) or sumr_134(5) or sumr_134(6) or sumr_134(7) or sumr_134(8));
E(376)<=not ( sumr_135(0) or sumr_135(1) or sumr_135(2) or sumr_135(3) or sumr_135(4) or sumr_135(5) or sumr_135(6) or sumr_135(7) or sumr_135(8));
E(375)<=not ( sumr_136(0) or sumr_136(1) or sumr_136(2) or sumr_136(3) or sumr_136(4) or sumr_136(5) or sumr_136(6) or sumr_136(7) or sumr_136(8));
E(374)<=not ( sumr_137(0) or sumr_137(1) or sumr_137(2) or sumr_137(3) or sumr_137(4) or sumr_137(5) or sumr_137(6) or sumr_137(7) or sumr_137(8));
E(373)<=not ( sumr_138(0) or sumr_138(1) or sumr_138(2) or sumr_138(3) or sumr_138(4) or sumr_138(5) or sumr_138(6) or sumr_138(7) or sumr_138(8));
E(372)<=not ( sumr_139(0) or sumr_139(1) or sumr_139(2) or sumr_139(3) or sumr_139(4) or sumr_139(5) or sumr_139(6) or sumr_139(7) or sumr_139(8));
E(371)<=not ( sumr_140(0) or sumr_140(1) or sumr_140(2) or sumr_140(3) or sumr_140(4) or sumr_140(5) or sumr_140(6) or sumr_140(7) or sumr_140(8));
E(370)<=not ( sumr_141(0) or sumr_141(1) or sumr_141(2) or sumr_141(3) or sumr_141(4) or sumr_141(5) or sumr_141(6) or sumr_141(7) or sumr_141(8));
E(369)<=not ( sumr_142(0) or sumr_142(1) or sumr_142(2) or sumr_142(3) or sumr_142(4) or sumr_142(5) or sumr_142(6) or sumr_142(7) or sumr_142(8));
E(368)<=not ( sumr_143(0) or sumr_143(1) or sumr_143(2) or sumr_143(3) or sumr_143(4) or sumr_143(5) or sumr_143(6) or sumr_143(7) or sumr_143(8));
E(367)<=not ( sumr_144(0) or sumr_144(1) or sumr_144(2) or sumr_144(3) or sumr_144(4) or sumr_144(5) or sumr_144(6) or sumr_144(7) or sumr_144(8));
E(366)<=not ( sumr_145(0) or sumr_145(1) or sumr_145(2) or sumr_145(3) or sumr_145(4) or sumr_145(5) or sumr_145(6) or sumr_145(7) or sumr_145(8));
E(365)<=not ( sumr_146(0) or sumr_146(1) or sumr_146(2) or sumr_146(3) or sumr_146(4) or sumr_146(5) or sumr_146(6) or sumr_146(7) or sumr_146(8));
E(364)<=not ( sumr_147(0) or sumr_147(1) or sumr_147(2) or sumr_147(3) or sumr_147(4) or sumr_147(5) or sumr_147(6) or sumr_147(7) or sumr_147(8));
E(363)<=not ( sumr_148(0) or sumr_148(1) or sumr_148(2) or sumr_148(3) or sumr_148(4) or sumr_148(5) or sumr_148(6) or sumr_148(7) or sumr_148(8));
E(362)<=not ( sumr_149(0) or sumr_149(1) or sumr_149(2) or sumr_149(3) or sumr_149(4) or sumr_149(5) or sumr_149(6) or sumr_149(7) or sumr_149(8));
E(361)<=not ( sumr_150(0) or sumr_150(1) or sumr_150(2) or sumr_150(3) or sumr_150(4) or sumr_150(5) or sumr_150(6) or sumr_150(7) or sumr_150(8));
E(360)<=not ( sumr_151(0) or sumr_151(1) or sumr_151(2) or sumr_151(3) or sumr_151(4) or sumr_151(5) or sumr_151(6) or sumr_151(7) or sumr_151(8));
E(359)<=not ( sumr_152(0) or sumr_152(1) or sumr_152(2) or sumr_152(3) or sumr_152(4) or sumr_152(5) or sumr_152(6) or sumr_152(7) or sumr_152(8));
E(358)<=not ( sumr_153(0) or sumr_153(1) or sumr_153(2) or sumr_153(3) or sumr_153(4) or sumr_153(5) or sumr_153(6) or sumr_153(7) or sumr_153(8));
E(357)<=not ( sumr_154(0) or sumr_154(1) or sumr_154(2) or sumr_154(3) or sumr_154(4) or sumr_154(5) or sumr_154(6) or sumr_154(7) or sumr_154(8));
E(356)<=not ( sumr_155(0) or sumr_155(1) or sumr_155(2) or sumr_155(3) or sumr_155(4) or sumr_155(5) or sumr_155(6) or sumr_155(7) or sumr_155(8));
E(355)<=not ( sumr_156(0) or sumr_156(1) or sumr_156(2) or sumr_156(3) or sumr_156(4) or sumr_156(5) or sumr_156(6) or sumr_156(7) or sumr_156(8));
E(354)<=not ( sumr_157(0) or sumr_157(1) or sumr_157(2) or sumr_157(3) or sumr_157(4) or sumr_157(5) or sumr_157(6) or sumr_157(7) or sumr_157(8));
E(353)<=not ( sumr_158(0) or sumr_158(1) or sumr_158(2) or sumr_158(3) or sumr_158(4) or sumr_158(5) or sumr_158(6) or sumr_158(7) or sumr_158(8));
E(352)<=not ( sumr_159(0) or sumr_159(1) or sumr_159(2) or sumr_159(3) or sumr_159(4) or sumr_159(5) or sumr_159(6) or sumr_159(7) or sumr_159(8));
E(351)<=not ( sumr_160(0) or sumr_160(1) or sumr_160(2) or sumr_160(3) or sumr_160(4) or sumr_160(5) or sumr_160(6) or sumr_160(7) or sumr_160(8));
E(350)<=not ( sumr_161(0) or sumr_161(1) or sumr_161(2) or sumr_161(3) or sumr_161(4) or sumr_161(5) or sumr_161(6) or sumr_161(7) or sumr_161(8));
E(349)<=not ( sumr_162(0) or sumr_162(1) or sumr_162(2) or sumr_162(3) or sumr_162(4) or sumr_162(5) or sumr_162(6) or sumr_162(7) or sumr_162(8));
E(348)<=not ( sumr_163(0) or sumr_163(1) or sumr_163(2) or sumr_163(3) or sumr_163(4) or sumr_163(5) or sumr_163(6) or sumr_163(7) or sumr_163(8));
E(347)<=not ( sumr_164(0) or sumr_164(1) or sumr_164(2) or sumr_164(3) or sumr_164(4) or sumr_164(5) or sumr_164(6) or sumr_164(7) or sumr_164(8));
E(346)<=not ( sumr_165(0) or sumr_165(1) or sumr_165(2) or sumr_165(3) or sumr_165(4) or sumr_165(5) or sumr_165(6) or sumr_165(7) or sumr_165(8));
E(345)<=not ( sumr_166(0) or sumr_166(1) or sumr_166(2) or sumr_166(3) or sumr_166(4) or sumr_166(5) or sumr_166(6) or sumr_166(7) or sumr_166(8));
E(344)<=not ( sumr_167(0) or sumr_167(1) or sumr_167(2) or sumr_167(3) or sumr_167(4) or sumr_167(5) or sumr_167(6) or sumr_167(7) or sumr_167(8));
E(343)<=not ( sumr_168(0) or sumr_168(1) or sumr_168(2) or sumr_168(3) or sumr_168(4) or sumr_168(5) or sumr_168(6) or sumr_168(7) or sumr_168(8));
E(342)<=not ( sumr_169(0) or sumr_169(1) or sumr_169(2) or sumr_169(3) or sumr_169(4) or sumr_169(5) or sumr_169(6) or sumr_169(7) or sumr_169(8));
E(341)<=not ( sumr_170(0) or sumr_170(1) or sumr_170(2) or sumr_170(3) or sumr_170(4) or sumr_170(5) or sumr_170(6) or sumr_170(7) or sumr_170(8));
E(340)<=not ( sumr_171(0) or sumr_171(1) or sumr_171(2) or sumr_171(3) or sumr_171(4) or sumr_171(5) or sumr_171(6) or sumr_171(7) or sumr_171(8));
E(339)<=not ( sumr_172(0) or sumr_172(1) or sumr_172(2) or sumr_172(3) or sumr_172(4) or sumr_172(5) or sumr_172(6) or sumr_172(7) or sumr_172(8));
E(338)<=not ( sumr_173(0) or sumr_173(1) or sumr_173(2) or sumr_173(3) or sumr_173(4) or sumr_173(5) or sumr_173(6) or sumr_173(7) or sumr_173(8));
E(337)<=not ( sumr_174(0) or sumr_174(1) or sumr_174(2) or sumr_174(3) or sumr_174(4) or sumr_174(5) or sumr_174(6) or sumr_174(7) or sumr_174(8));
E(336)<=not ( sumr_175(0) or sumr_175(1) or sumr_175(2) or sumr_175(3) or sumr_175(4) or sumr_175(5) or sumr_175(6) or sumr_175(7) or sumr_175(8));
E(335)<=not ( sumr_176(0) or sumr_176(1) or sumr_176(2) or sumr_176(3) or sumr_176(4) or sumr_176(5) or sumr_176(6) or sumr_176(7) or sumr_176(8));
E(334)<=not ( sumr_177(0) or sumr_177(1) or sumr_177(2) or sumr_177(3) or sumr_177(4) or sumr_177(5) or sumr_177(6) or sumr_177(7) or sumr_177(8));
E(333)<=not ( sumr_178(0) or sumr_178(1) or sumr_178(2) or sumr_178(3) or sumr_178(4) or sumr_178(5) or sumr_178(6) or sumr_178(7) or sumr_178(8));
E(332)<=not ( sumr_179(0) or sumr_179(1) or sumr_179(2) or sumr_179(3) or sumr_179(4) or sumr_179(5) or sumr_179(6) or sumr_179(7) or sumr_179(8));
E(331)<=not ( sumr_180(0) or sumr_180(1) or sumr_180(2) or sumr_180(3) or sumr_180(4) or sumr_180(5) or sumr_180(6) or sumr_180(7) or sumr_180(8));
E(330)<=not ( sumr_181(0) or sumr_181(1) or sumr_181(2) or sumr_181(3) or sumr_181(4) or sumr_181(5) or sumr_181(6) or sumr_181(7) or sumr_181(8));
E(329)<=not ( sumr_182(0) or sumr_182(1) or sumr_182(2) or sumr_182(3) or sumr_182(4) or sumr_182(5) or sumr_182(6) or sumr_182(7) or sumr_182(8));
E(328)<=not ( sumr_183(0) or sumr_183(1) or sumr_183(2) or sumr_183(3) or sumr_183(4) or sumr_183(5) or sumr_183(6) or sumr_183(7) or sumr_183(8));
E(327)<=not ( sumr_184(0) or sumr_184(1) or sumr_184(2) or sumr_184(3) or sumr_184(4) or sumr_184(5) or sumr_184(6) or sumr_184(7) or sumr_184(8));
E(326)<=not ( sumr_185(0) or sumr_185(1) or sumr_185(2) or sumr_185(3) or sumr_185(4) or sumr_185(5) or sumr_185(6) or sumr_185(7) or sumr_185(8));
E(325)<=not ( sumr_186(0) or sumr_186(1) or sumr_186(2) or sumr_186(3) or sumr_186(4) or sumr_186(5) or sumr_186(6) or sumr_186(7) or sumr_186(8));
E(324)<=not ( sumr_187(0) or sumr_187(1) or sumr_187(2) or sumr_187(3) or sumr_187(4) or sumr_187(5) or sumr_187(6) or sumr_187(7) or sumr_187(8));
E(323)<=not ( sumr_188(0) or sumr_188(1) or sumr_188(2) or sumr_188(3) or sumr_188(4) or sumr_188(5) or sumr_188(6) or sumr_188(7) or sumr_188(8));
E(322)<=not ( sumr_189(0) or sumr_189(1) or sumr_189(2) or sumr_189(3) or sumr_189(4) or sumr_189(5) or sumr_189(6) or sumr_189(7) or sumr_189(8));
E(321)<=not ( sumr_190(0) or sumr_190(1) or sumr_190(2) or sumr_190(3) or sumr_190(4) or sumr_190(5) or sumr_190(6) or sumr_190(7) or sumr_190(8));
E(320)<=not ( sumr_191(0) or sumr_191(1) or sumr_191(2) or sumr_191(3) or sumr_191(4) or sumr_191(5) or sumr_191(6) or sumr_191(7) or sumr_191(8));
E(319)<=not ( sumr_192(0) or sumr_192(1) or sumr_192(2) or sumr_192(3) or sumr_192(4) or sumr_192(5) or sumr_192(6) or sumr_192(7) or sumr_192(8));
E(318)<=not ( sumr_193(0) or sumr_193(1) or sumr_193(2) or sumr_193(3) or sumr_193(4) or sumr_193(5) or sumr_193(6) or sumr_193(7) or sumr_193(8));
E(317)<=not ( sumr_194(0) or sumr_194(1) or sumr_194(2) or sumr_194(3) or sumr_194(4) or sumr_194(5) or sumr_194(6) or sumr_194(7) or sumr_194(8));
E(316)<=not ( sumr_195(0) or sumr_195(1) or sumr_195(2) or sumr_195(3) or sumr_195(4) or sumr_195(5) or sumr_195(6) or sumr_195(7) or sumr_195(8));
E(315)<=not ( sumr_196(0) or sumr_196(1) or sumr_196(2) or sumr_196(3) or sumr_196(4) or sumr_196(5) or sumr_196(6) or sumr_196(7) or sumr_196(8));
E(314)<=not ( sumr_197(0) or sumr_197(1) or sumr_197(2) or sumr_197(3) or sumr_197(4) or sumr_197(5) or sumr_197(6) or sumr_197(7) or sumr_197(8));
E(313)<=not ( sumr_198(0) or sumr_198(1) or sumr_198(2) or sumr_198(3) or sumr_198(4) or sumr_198(5) or sumr_198(6) or sumr_198(7) or sumr_198(8));
E(312)<=not ( sumr_199(0) or sumr_199(1) or sumr_199(2) or sumr_199(3) or sumr_199(4) or sumr_199(5) or sumr_199(6) or sumr_199(7) or sumr_199(8));
E(311)<=not ( sumr_200(0) or sumr_200(1) or sumr_200(2) or sumr_200(3) or sumr_200(4) or sumr_200(5) or sumr_200(6) or sumr_200(7) or sumr_200(8));
E(310)<=not ( sumr_201(0) or sumr_201(1) or sumr_201(2) or sumr_201(3) or sumr_201(4) or sumr_201(5) or sumr_201(6) or sumr_201(7) or sumr_201(8));
E(309)<=not ( sumr_202(0) or sumr_202(1) or sumr_202(2) or sumr_202(3) or sumr_202(4) or sumr_202(5) or sumr_202(6) or sumr_202(7) or sumr_202(8));
E(308)<=not ( sumr_203(0) or sumr_203(1) or sumr_203(2) or sumr_203(3) or sumr_203(4) or sumr_203(5) or sumr_203(6) or sumr_203(7) or sumr_203(8));
E(307)<=not ( sumr_204(0) or sumr_204(1) or sumr_204(2) or sumr_204(3) or sumr_204(4) or sumr_204(5) or sumr_204(6) or sumr_204(7) or sumr_204(8));
E(306)<=not ( sumr_205(0) or sumr_205(1) or sumr_205(2) or sumr_205(3) or sumr_205(4) or sumr_205(5) or sumr_205(6) or sumr_205(7) or sumr_205(8));
E(305)<=not ( sumr_206(0) or sumr_206(1) or sumr_206(2) or sumr_206(3) or sumr_206(4) or sumr_206(5) or sumr_206(6) or sumr_206(7) or sumr_206(8));
E(304)<=not ( sumr_207(0) or sumr_207(1) or sumr_207(2) or sumr_207(3) or sumr_207(4) or sumr_207(5) or sumr_207(6) or sumr_207(7) or sumr_207(8));
E(303)<=not ( sumr_208(0) or sumr_208(1) or sumr_208(2) or sumr_208(3) or sumr_208(4) or sumr_208(5) or sumr_208(6) or sumr_208(7) or sumr_208(8));
E(302)<=not ( sumr_209(0) or sumr_209(1) or sumr_209(2) or sumr_209(3) or sumr_209(4) or sumr_209(5) or sumr_209(6) or sumr_209(7) or sumr_209(8));
E(301)<=not ( sumr_210(0) or sumr_210(1) or sumr_210(2) or sumr_210(3) or sumr_210(4) or sumr_210(5) or sumr_210(6) or sumr_210(7) or sumr_210(8));
E(300)<=not ( sumr_211(0) or sumr_211(1) or sumr_211(2) or sumr_211(3) or sumr_211(4) or sumr_211(5) or sumr_211(6) or sumr_211(7) or sumr_211(8));
E(299)<=not ( sumr_212(0) or sumr_212(1) or sumr_212(2) or sumr_212(3) or sumr_212(4) or sumr_212(5) or sumr_212(6) or sumr_212(7) or sumr_212(8));
E(298)<=not ( sumr_213(0) or sumr_213(1) or sumr_213(2) or sumr_213(3) or sumr_213(4) or sumr_213(5) or sumr_213(6) or sumr_213(7) or sumr_213(8));
E(297)<=not ( sumr_214(0) or sumr_214(1) or sumr_214(2) or sumr_214(3) or sumr_214(4) or sumr_214(5) or sumr_214(6) or sumr_214(7) or sumr_214(8));
E(296)<=not ( sumr_215(0) or sumr_215(1) or sumr_215(2) or sumr_215(3) or sumr_215(4) or sumr_215(5) or sumr_215(6) or sumr_215(7) or sumr_215(8));
E(295)<=not ( sumr_216(0) or sumr_216(1) or sumr_216(2) or sumr_216(3) or sumr_216(4) or sumr_216(5) or sumr_216(6) or sumr_216(7) or sumr_216(8));
E(294)<=not ( sumr_217(0) or sumr_217(1) or sumr_217(2) or sumr_217(3) or sumr_217(4) or sumr_217(5) or sumr_217(6) or sumr_217(7) or sumr_217(8));
E(293)<=not ( sumr_218(0) or sumr_218(1) or sumr_218(2) or sumr_218(3) or sumr_218(4) or sumr_218(5) or sumr_218(6) or sumr_218(7) or sumr_218(8));
E(292)<=not ( sumr_219(0) or sumr_219(1) or sumr_219(2) or sumr_219(3) or sumr_219(4) or sumr_219(5) or sumr_219(6) or sumr_219(7) or sumr_219(8));
E(291)<=not ( sumr_220(0) or sumr_220(1) or sumr_220(2) or sumr_220(3) or sumr_220(4) or sumr_220(5) or sumr_220(6) or sumr_220(7) or sumr_220(8));
E(290)<=not ( sumr_221(0) or sumr_221(1) or sumr_221(2) or sumr_221(3) or sumr_221(4) or sumr_221(5) or sumr_221(6) or sumr_221(7) or sumr_221(8));
E(289)<=not ( sumr_222(0) or sumr_222(1) or sumr_222(2) or sumr_222(3) or sumr_222(4) or sumr_222(5) or sumr_222(6) or sumr_222(7) or sumr_222(8));
E(288)<=not ( sumr_223(0) or sumr_223(1) or sumr_223(2) or sumr_223(3) or sumr_223(4) or sumr_223(5) or sumr_223(6) or sumr_223(7) or sumr_223(8));
E(287)<=not ( sumr_224(0) or sumr_224(1) or sumr_224(2) or sumr_224(3) or sumr_224(4) or sumr_224(5) or sumr_224(6) or sumr_224(7) or sumr_224(8));
E(286)<=not ( sumr_225(0) or sumr_225(1) or sumr_225(2) or sumr_225(3) or sumr_225(4) or sumr_225(5) or sumr_225(6) or sumr_225(7) or sumr_225(8));
E(285)<=not ( sumr_226(0) or sumr_226(1) or sumr_226(2) or sumr_226(3) or sumr_226(4) or sumr_226(5) or sumr_226(6) or sumr_226(7) or sumr_226(8));
E(284)<=not ( sumr_227(0) or sumr_227(1) or sumr_227(2) or sumr_227(3) or sumr_227(4) or sumr_227(5) or sumr_227(6) or sumr_227(7) or sumr_227(8));
E(283)<=not ( sumr_228(0) or sumr_228(1) or sumr_228(2) or sumr_228(3) or sumr_228(4) or sumr_228(5) or sumr_228(6) or sumr_228(7) or sumr_228(8));
E(282)<=not ( sumr_229(0) or sumr_229(1) or sumr_229(2) or sumr_229(3) or sumr_229(4) or sumr_229(5) or sumr_229(6) or sumr_229(7) or sumr_229(8));
E(281)<=not ( sumr_230(0) or sumr_230(1) or sumr_230(2) or sumr_230(3) or sumr_230(4) or sumr_230(5) or sumr_230(6) or sumr_230(7) or sumr_230(8));
E(280)<=not ( sumr_231(0) or sumr_231(1) or sumr_231(2) or sumr_231(3) or sumr_231(4) or sumr_231(5) or sumr_231(6) or sumr_231(7) or sumr_231(8));
E(279)<=not ( sumr_232(0) or sumr_232(1) or sumr_232(2) or sumr_232(3) or sumr_232(4) or sumr_232(5) or sumr_232(6) or sumr_232(7) or sumr_232(8));
E(278)<=not ( sumr_233(0) or sumr_233(1) or sumr_233(2) or sumr_233(3) or sumr_233(4) or sumr_233(5) or sumr_233(6) or sumr_233(7) or sumr_233(8));
E(277)<=not ( sumr_234(0) or sumr_234(1) or sumr_234(2) or sumr_234(3) or sumr_234(4) or sumr_234(5) or sumr_234(6) or sumr_234(7) or sumr_234(8));
E(276)<=not ( sumr_235(0) or sumr_235(1) or sumr_235(2) or sumr_235(3) or sumr_235(4) or sumr_235(5) or sumr_235(6) or sumr_235(7) or sumr_235(8));
E(275)<=not ( sumr_236(0) or sumr_236(1) or sumr_236(2) or sumr_236(3) or sumr_236(4) or sumr_236(5) or sumr_236(6) or sumr_236(7) or sumr_236(8));
E(274)<=not ( sumr_237(0) or sumr_237(1) or sumr_237(2) or sumr_237(3) or sumr_237(4) or sumr_237(5) or sumr_237(6) or sumr_237(7) or sumr_237(8));
E(273)<=not ( sumr_238(0) or sumr_238(1) or sumr_238(2) or sumr_238(3) or sumr_238(4) or sumr_238(5) or sumr_238(6) or sumr_238(7) or sumr_238(8));
E(272)<=not ( sumr_239(0) or sumr_239(1) or sumr_239(2) or sumr_239(3) or sumr_239(4) or sumr_239(5) or sumr_239(6) or sumr_239(7) or sumr_239(8));
E(271)<=not ( sumr_240(0) or sumr_240(1) or sumr_240(2) or sumr_240(3) or sumr_240(4) or sumr_240(5) or sumr_240(6) or sumr_240(7) or sumr_240(8));
E(270)<=not ( sumr_241(0) or sumr_241(1) or sumr_241(2) or sumr_241(3) or sumr_241(4) or sumr_241(5) or sumr_241(6) or sumr_241(7) or sumr_241(8));
E(269)<=not ( sumr_242(0) or sumr_242(1) or sumr_242(2) or sumr_242(3) or sumr_242(4) or sumr_242(5) or sumr_242(6) or sumr_242(7) or sumr_242(8));
E(268)<=not ( sumr_243(0) or sumr_243(1) or sumr_243(2) or sumr_243(3) or sumr_243(4) or sumr_243(5) or sumr_243(6) or sumr_243(7) or sumr_243(8));
E(267)<=not ( sumr_244(0) or sumr_244(1) or sumr_244(2) or sumr_244(3) or sumr_244(4) or sumr_244(5) or sumr_244(6) or sumr_244(7) or sumr_244(8));
E(266)<=not ( sumr_245(0) or sumr_245(1) or sumr_245(2) or sumr_245(3) or sumr_245(4) or sumr_245(5) or sumr_245(6) or sumr_245(7) or sumr_245(8));
E(265)<=not ( sumr_246(0) or sumr_246(1) or sumr_246(2) or sumr_246(3) or sumr_246(4) or sumr_246(5) or sumr_246(6) or sumr_246(7) or sumr_246(8));
E(264)<=not ( sumr_247(0) or sumr_247(1) or sumr_247(2) or sumr_247(3) or sumr_247(4) or sumr_247(5) or sumr_247(6) or sumr_247(7) or sumr_247(8));
E(263)<=not ( sumr_248(0) or sumr_248(1) or sumr_248(2) or sumr_248(3) or sumr_248(4) or sumr_248(5) or sumr_248(6) or sumr_248(7) or sumr_248(8));
E(262)<=not ( sumr_249(0) or sumr_249(1) or sumr_249(2) or sumr_249(3) or sumr_249(4) or sumr_249(5) or sumr_249(6) or sumr_249(7) or sumr_249(8));
E(261)<=not ( sumr_250(0) or sumr_250(1) or sumr_250(2) or sumr_250(3) or sumr_250(4) or sumr_250(5) or sumr_250(6) or sumr_250(7) or sumr_250(8));
E(260)<=not ( sumr_251(0) or sumr_251(1) or sumr_251(2) or sumr_251(3) or sumr_251(4) or sumr_251(5) or sumr_251(6) or sumr_251(7) or sumr_251(8));
E(259)<=not ( sumr_252(0) or sumr_252(1) or sumr_252(2) or sumr_252(3) or sumr_252(4) or sumr_252(5) or sumr_252(6) or sumr_252(7) or sumr_252(8));
E(258)<=not ( sumr_253(0) or sumr_253(1) or sumr_253(2) or sumr_253(3) or sumr_253(4) or sumr_253(5) or sumr_253(6) or sumr_253(7) or sumr_253(8));
E(257)<=not ( sumr_254(0) or sumr_254(1) or sumr_254(2) or sumr_254(3) or sumr_254(4) or sumr_254(5) or sumr_254(6) or sumr_254(7) or sumr_254(8));
E(256)<=not ( sumr_255(0) or sumr_255(1) or sumr_255(2) or sumr_255(3) or sumr_255(4) or sumr_255(5) or sumr_255(6) or sumr_255(7) or sumr_255(8));
E(255)<=not ( sumr_256(0) or sumr_256(1) or sumr_256(2) or sumr_256(3) or sumr_256(4) or sumr_256(5) or sumr_256(6) or sumr_256(7) or sumr_256(8));
E(254)<=not ( sumr_257(0) or sumr_257(1) or sumr_257(2) or sumr_257(3) or sumr_257(4) or sumr_257(5) or sumr_257(6) or sumr_257(7) or sumr_257(8));
E(253)<=not ( sumr_258(0) or sumr_258(1) or sumr_258(2) or sumr_258(3) or sumr_258(4) or sumr_258(5) or sumr_258(6) or sumr_258(7) or sumr_258(8));
E(252)<=not ( sumr_259(0) or sumr_259(1) or sumr_259(2) or sumr_259(3) or sumr_259(4) or sumr_259(5) or sumr_259(6) or sumr_259(7) or sumr_259(8));
E(251)<=not ( sumr_260(0) or sumr_260(1) or sumr_260(2) or sumr_260(3) or sumr_260(4) or sumr_260(5) or sumr_260(6) or sumr_260(7) or sumr_260(8));
E(250)<=not ( sumr_261(0) or sumr_261(1) or sumr_261(2) or sumr_261(3) or sumr_261(4) or sumr_261(5) or sumr_261(6) or sumr_261(7) or sumr_261(8));
E(249)<=not ( sumr_262(0) or sumr_262(1) or sumr_262(2) or sumr_262(3) or sumr_262(4) or sumr_262(5) or sumr_262(6) or sumr_262(7) or sumr_262(8));
E(248)<=not ( sumr_263(0) or sumr_263(1) or sumr_263(2) or sumr_263(3) or sumr_263(4) or sumr_263(5) or sumr_263(6) or sumr_263(7) or sumr_263(8));
E(247)<=not ( sumr_264(0) or sumr_264(1) or sumr_264(2) or sumr_264(3) or sumr_264(4) or sumr_264(5) or sumr_264(6) or sumr_264(7) or sumr_264(8));
E(246)<=not ( sumr_265(0) or sumr_265(1) or sumr_265(2) or sumr_265(3) or sumr_265(4) or sumr_265(5) or sumr_265(6) or sumr_265(7) or sumr_265(8));
E(245)<=not ( sumr_266(0) or sumr_266(1) or sumr_266(2) or sumr_266(3) or sumr_266(4) or sumr_266(5) or sumr_266(6) or sumr_266(7) or sumr_266(8));
E(244)<=not ( sumr_267(0) or sumr_267(1) or sumr_267(2) or sumr_267(3) or sumr_267(4) or sumr_267(5) or sumr_267(6) or sumr_267(7) or sumr_267(8));
E(243)<=not ( sumr_268(0) or sumr_268(1) or sumr_268(2) or sumr_268(3) or sumr_268(4) or sumr_268(5) or sumr_268(6) or sumr_268(7) or sumr_268(8));
E(242)<=not ( sumr_269(0) or sumr_269(1) or sumr_269(2) or sumr_269(3) or sumr_269(4) or sumr_269(5) or sumr_269(6) or sumr_269(7) or sumr_269(8));
E(241)<=not ( sumr_270(0) or sumr_270(1) or sumr_270(2) or sumr_270(3) or sumr_270(4) or sumr_270(5) or sumr_270(6) or sumr_270(7) or sumr_270(8));
E(240)<=not ( sumr_271(0) or sumr_271(1) or sumr_271(2) or sumr_271(3) or sumr_271(4) or sumr_271(5) or sumr_271(6) or sumr_271(7) or sumr_271(8));
E(239)<=not ( sumr_272(0) or sumr_272(1) or sumr_272(2) or sumr_272(3) or sumr_272(4) or sumr_272(5) or sumr_272(6) or sumr_272(7) or sumr_272(8));
E(238)<=not ( sumr_273(0) or sumr_273(1) or sumr_273(2) or sumr_273(3) or sumr_273(4) or sumr_273(5) or sumr_273(6) or sumr_273(7) or sumr_273(8));
E(237)<=not ( sumr_274(0) or sumr_274(1) or sumr_274(2) or sumr_274(3) or sumr_274(4) or sumr_274(5) or sumr_274(6) or sumr_274(7) or sumr_274(8));
E(236)<=not ( sumr_275(0) or sumr_275(1) or sumr_275(2) or sumr_275(3) or sumr_275(4) or sumr_275(5) or sumr_275(6) or sumr_275(7) or sumr_275(8));
E(235)<=not ( sumr_276(0) or sumr_276(1) or sumr_276(2) or sumr_276(3) or sumr_276(4) or sumr_276(5) or sumr_276(6) or sumr_276(7) or sumr_276(8));
E(234)<=not ( sumr_277(0) or sumr_277(1) or sumr_277(2) or sumr_277(3) or sumr_277(4) or sumr_277(5) or sumr_277(6) or sumr_277(7) or sumr_277(8));
E(233)<=not ( sumr_278(0) or sumr_278(1) or sumr_278(2) or sumr_278(3) or sumr_278(4) or sumr_278(5) or sumr_278(6) or sumr_278(7) or sumr_278(8));
E(232)<=not ( sumr_279(0) or sumr_279(1) or sumr_279(2) or sumr_279(3) or sumr_279(4) or sumr_279(5) or sumr_279(6) or sumr_279(7) or sumr_279(8));
E(231)<=not ( sumr_280(0) or sumr_280(1) or sumr_280(2) or sumr_280(3) or sumr_280(4) or sumr_280(5) or sumr_280(6) or sumr_280(7) or sumr_280(8));
E(230)<=not ( sumr_281(0) or sumr_281(1) or sumr_281(2) or sumr_281(3) or sumr_281(4) or sumr_281(5) or sumr_281(6) or sumr_281(7) or sumr_281(8));
E(229)<=not ( sumr_282(0) or sumr_282(1) or sumr_282(2) or sumr_282(3) or sumr_282(4) or sumr_282(5) or sumr_282(6) or sumr_282(7) or sumr_282(8));
E(228)<=not ( sumr_283(0) or sumr_283(1) or sumr_283(2) or sumr_283(3) or sumr_283(4) or sumr_283(5) or sumr_283(6) or sumr_283(7) or sumr_283(8));
E(227)<=not ( sumr_284(0) or sumr_284(1) or sumr_284(2) or sumr_284(3) or sumr_284(4) or sumr_284(5) or sumr_284(6) or sumr_284(7) or sumr_284(8));
E(226)<=not ( sumr_285(0) or sumr_285(1) or sumr_285(2) or sumr_285(3) or sumr_285(4) or sumr_285(5) or sumr_285(6) or sumr_285(7) or sumr_285(8));
E(225)<=not ( sumr_286(0) or sumr_286(1) or sumr_286(2) or sumr_286(3) or sumr_286(4) or sumr_286(5) or sumr_286(6) or sumr_286(7) or sumr_286(8));
E(224)<=not ( sumr_287(0) or sumr_287(1) or sumr_287(2) or sumr_287(3) or sumr_287(4) or sumr_287(5) or sumr_287(6) or sumr_287(7) or sumr_287(8));
E(223)<=not ( sumr_288(0) or sumr_288(1) or sumr_288(2) or sumr_288(3) or sumr_288(4) or sumr_288(5) or sumr_288(6) or sumr_288(7) or sumr_288(8));
E(222)<=not ( sumr_289(0) or sumr_289(1) or sumr_289(2) or sumr_289(3) or sumr_289(4) or sumr_289(5) or sumr_289(6) or sumr_289(7) or sumr_289(8));
E(221)<=not ( sumr_290(0) or sumr_290(1) or sumr_290(2) or sumr_290(3) or sumr_290(4) or sumr_290(5) or sumr_290(6) or sumr_290(7) or sumr_290(8));
E(220)<=not ( sumr_291(0) or sumr_291(1) or sumr_291(2) or sumr_291(3) or sumr_291(4) or sumr_291(5) or sumr_291(6) or sumr_291(7) or sumr_291(8));
E(219)<=not ( sumr_292(0) or sumr_292(1) or sumr_292(2) or sumr_292(3) or sumr_292(4) or sumr_292(5) or sumr_292(6) or sumr_292(7) or sumr_292(8));
E(218)<=not ( sumr_293(0) or sumr_293(1) or sumr_293(2) or sumr_293(3) or sumr_293(4) or sumr_293(5) or sumr_293(6) or sumr_293(7) or sumr_293(8));
E(217)<=not ( sumr_294(0) or sumr_294(1) or sumr_294(2) or sumr_294(3) or sumr_294(4) or sumr_294(5) or sumr_294(6) or sumr_294(7) or sumr_294(8));
E(216)<=not ( sumr_295(0) or sumr_295(1) or sumr_295(2) or sumr_295(3) or sumr_295(4) or sumr_295(5) or sumr_295(6) or sumr_295(7) or sumr_295(8));
E(215)<=not ( sumr_296(0) or sumr_296(1) or sumr_296(2) or sumr_296(3) or sumr_296(4) or sumr_296(5) or sumr_296(6) or sumr_296(7) or sumr_296(8));
E(214)<=not ( sumr_297(0) or sumr_297(1) or sumr_297(2) or sumr_297(3) or sumr_297(4) or sumr_297(5) or sumr_297(6) or sumr_297(7) or sumr_297(8));
E(213)<=not ( sumr_298(0) or sumr_298(1) or sumr_298(2) or sumr_298(3) or sumr_298(4) or sumr_298(5) or sumr_298(6) or sumr_298(7) or sumr_298(8));
E(212)<=not ( sumr_299(0) or sumr_299(1) or sumr_299(2) or sumr_299(3) or sumr_299(4) or sumr_299(5) or sumr_299(6) or sumr_299(7) or sumr_299(8));
E(211)<=not ( sumr_300(0) or sumr_300(1) or sumr_300(2) or sumr_300(3) or sumr_300(4) or sumr_300(5) or sumr_300(6) or sumr_300(7) or sumr_300(8));
E(210)<=not ( sumr_301(0) or sumr_301(1) or sumr_301(2) or sumr_301(3) or sumr_301(4) or sumr_301(5) or sumr_301(6) or sumr_301(7) or sumr_301(8));
E(209)<=not ( sumr_302(0) or sumr_302(1) or sumr_302(2) or sumr_302(3) or sumr_302(4) or sumr_302(5) or sumr_302(6) or sumr_302(7) or sumr_302(8));
E(208)<=not ( sumr_303(0) or sumr_303(1) or sumr_303(2) or sumr_303(3) or sumr_303(4) or sumr_303(5) or sumr_303(6) or sumr_303(7) or sumr_303(8));
E(207)<=not ( sumr_304(0) or sumr_304(1) or sumr_304(2) or sumr_304(3) or sumr_304(4) or sumr_304(5) or sumr_304(6) or sumr_304(7) or sumr_304(8));
E(206)<=not ( sumr_305(0) or sumr_305(1) or sumr_305(2) or sumr_305(3) or sumr_305(4) or sumr_305(5) or sumr_305(6) or sumr_305(7) or sumr_305(8));
E(205)<=not ( sumr_306(0) or sumr_306(1) or sumr_306(2) or sumr_306(3) or sumr_306(4) or sumr_306(5) or sumr_306(6) or sumr_306(7) or sumr_306(8));
E(204)<=not ( sumr_307(0) or sumr_307(1) or sumr_307(2) or sumr_307(3) or sumr_307(4) or sumr_307(5) or sumr_307(6) or sumr_307(7) or sumr_307(8));
E(203)<=not ( sumr_308(0) or sumr_308(1) or sumr_308(2) or sumr_308(3) or sumr_308(4) or sumr_308(5) or sumr_308(6) or sumr_308(7) or sumr_308(8));
E(202)<=not ( sumr_309(0) or sumr_309(1) or sumr_309(2) or sumr_309(3) or sumr_309(4) or sumr_309(5) or sumr_309(6) or sumr_309(7) or sumr_309(8));
E(201)<=not ( sumr_310(0) or sumr_310(1) or sumr_310(2) or sumr_310(3) or sumr_310(4) or sumr_310(5) or sumr_310(6) or sumr_310(7) or sumr_310(8));
E(200)<=not ( sumr_311(0) or sumr_311(1) or sumr_311(2) or sumr_311(3) or sumr_311(4) or sumr_311(5) or sumr_311(6) or sumr_311(7) or sumr_311(8));
E(199)<=not ( sumr_312(0) or sumr_312(1) or sumr_312(2) or sumr_312(3) or sumr_312(4) or sumr_312(5) or sumr_312(6) or sumr_312(7) or sumr_312(8));
E(198)<=not ( sumr_313(0) or sumr_313(1) or sumr_313(2) or sumr_313(3) or sumr_313(4) or sumr_313(5) or sumr_313(6) or sumr_313(7) or sumr_313(8));
E(197)<=not ( sumr_314(0) or sumr_314(1) or sumr_314(2) or sumr_314(3) or sumr_314(4) or sumr_314(5) or sumr_314(6) or sumr_314(7) or sumr_314(8));
E(196)<=not ( sumr_315(0) or sumr_315(1) or sumr_315(2) or sumr_315(3) or sumr_315(4) or sumr_315(5) or sumr_315(6) or sumr_315(7) or sumr_315(8));
E(195)<=not ( sumr_316(0) or sumr_316(1) or sumr_316(2) or sumr_316(3) or sumr_316(4) or sumr_316(5) or sumr_316(6) or sumr_316(7) or sumr_316(8));
E(194)<=not ( sumr_317(0) or sumr_317(1) or sumr_317(2) or sumr_317(3) or sumr_317(4) or sumr_317(5) or sumr_317(6) or sumr_317(7) or sumr_317(8));
E(193)<=not ( sumr_318(0) or sumr_318(1) or sumr_318(2) or sumr_318(3) or sumr_318(4) or sumr_318(5) or sumr_318(6) or sumr_318(7) or sumr_318(8));
E(192)<=not ( sumr_319(0) or sumr_319(1) or sumr_319(2) or sumr_319(3) or sumr_319(4) or sumr_319(5) or sumr_319(6) or sumr_319(7) or sumr_319(8));
E(191)<=not ( sumr_320(0) or sumr_320(1) or sumr_320(2) or sumr_320(3) or sumr_320(4) or sumr_320(5) or sumr_320(6) or sumr_320(7) or sumr_320(8));
E(190)<=not ( sumr_321(0) or sumr_321(1) or sumr_321(2) or sumr_321(3) or sumr_321(4) or sumr_321(5) or sumr_321(6) or sumr_321(7) or sumr_321(8));
E(189)<=not ( sumr_322(0) or sumr_322(1) or sumr_322(2) or sumr_322(3) or sumr_322(4) or sumr_322(5) or sumr_322(6) or sumr_322(7) or sumr_322(8));
E(188)<=not ( sumr_323(0) or sumr_323(1) or sumr_323(2) or sumr_323(3) or sumr_323(4) or sumr_323(5) or sumr_323(6) or sumr_323(7) or sumr_323(8));
E(187)<=not ( sumr_324(0) or sumr_324(1) or sumr_324(2) or sumr_324(3) or sumr_324(4) or sumr_324(5) or sumr_324(6) or sumr_324(7) or sumr_324(8));
E(186)<=not ( sumr_325(0) or sumr_325(1) or sumr_325(2) or sumr_325(3) or sumr_325(4) or sumr_325(5) or sumr_325(6) or sumr_325(7) or sumr_325(8));
E(185)<=not ( sumr_326(0) or sumr_326(1) or sumr_326(2) or sumr_326(3) or sumr_326(4) or sumr_326(5) or sumr_326(6) or sumr_326(7) or sumr_326(8));
E(184)<=not ( sumr_327(0) or sumr_327(1) or sumr_327(2) or sumr_327(3) or sumr_327(4) or sumr_327(5) or sumr_327(6) or sumr_327(7) or sumr_327(8));
E(183)<=not ( sumr_328(0) or sumr_328(1) or sumr_328(2) or sumr_328(3) or sumr_328(4) or sumr_328(5) or sumr_328(6) or sumr_328(7) or sumr_328(8));
E(182)<=not ( sumr_329(0) or sumr_329(1) or sumr_329(2) or sumr_329(3) or sumr_329(4) or sumr_329(5) or sumr_329(6) or sumr_329(7) or sumr_329(8));
E(181)<=not ( sumr_330(0) or sumr_330(1) or sumr_330(2) or sumr_330(3) or sumr_330(4) or sumr_330(5) or sumr_330(6) or sumr_330(7) or sumr_330(8));
E(180)<=not ( sumr_331(0) or sumr_331(1) or sumr_331(2) or sumr_331(3) or sumr_331(4) or sumr_331(5) or sumr_331(6) or sumr_331(7) or sumr_331(8));
E(179)<=not ( sumr_332(0) or sumr_332(1) or sumr_332(2) or sumr_332(3) or sumr_332(4) or sumr_332(5) or sumr_332(6) or sumr_332(7) or sumr_332(8));
E(178)<=not ( sumr_333(0) or sumr_333(1) or sumr_333(2) or sumr_333(3) or sumr_333(4) or sumr_333(5) or sumr_333(6) or sumr_333(7) or sumr_333(8));
E(177)<=not ( sumr_334(0) or sumr_334(1) or sumr_334(2) or sumr_334(3) or sumr_334(4) or sumr_334(5) or sumr_334(6) or sumr_334(7) or sumr_334(8));
E(176)<=not ( sumr_335(0) or sumr_335(1) or sumr_335(2) or sumr_335(3) or sumr_335(4) or sumr_335(5) or sumr_335(6) or sumr_335(7) or sumr_335(8));
E(175)<=not ( sumr_336(0) or sumr_336(1) or sumr_336(2) or sumr_336(3) or sumr_336(4) or sumr_336(5) or sumr_336(6) or sumr_336(7) or sumr_336(8));
E(174)<=not ( sumr_337(0) or sumr_337(1) or sumr_337(2) or sumr_337(3) or sumr_337(4) or sumr_337(5) or sumr_337(6) or sumr_337(7) or sumr_337(8));
E(173)<=not ( sumr_338(0) or sumr_338(1) or sumr_338(2) or sumr_338(3) or sumr_338(4) or sumr_338(5) or sumr_338(6) or sumr_338(7) or sumr_338(8));
E(172)<=not ( sumr_339(0) or sumr_339(1) or sumr_339(2) or sumr_339(3) or sumr_339(4) or sumr_339(5) or sumr_339(6) or sumr_339(7) or sumr_339(8));
E(171)<=not ( sumr_340(0) or sumr_340(1) or sumr_340(2) or sumr_340(3) or sumr_340(4) or sumr_340(5) or sumr_340(6) or sumr_340(7) or sumr_340(8));
E(170)<=not ( sumr_341(0) or sumr_341(1) or sumr_341(2) or sumr_341(3) or sumr_341(4) or sumr_341(5) or sumr_341(6) or sumr_341(7) or sumr_341(8));
E(169)<=not ( sumr_342(0) or sumr_342(1) or sumr_342(2) or sumr_342(3) or sumr_342(4) or sumr_342(5) or sumr_342(6) or sumr_342(7) or sumr_342(8));
E(168)<=not ( sumr_343(0) or sumr_343(1) or sumr_343(2) or sumr_343(3) or sumr_343(4) or sumr_343(5) or sumr_343(6) or sumr_343(7) or sumr_343(8));
E(167)<=not ( sumr_344(0) or sumr_344(1) or sumr_344(2) or sumr_344(3) or sumr_344(4) or sumr_344(5) or sumr_344(6) or sumr_344(7) or sumr_344(8));
E(166)<=not ( sumr_345(0) or sumr_345(1) or sumr_345(2) or sumr_345(3) or sumr_345(4) or sumr_345(5) or sumr_345(6) or sumr_345(7) or sumr_345(8));
E(165)<=not ( sumr_346(0) or sumr_346(1) or sumr_346(2) or sumr_346(3) or sumr_346(4) or sumr_346(5) or sumr_346(6) or sumr_346(7) or sumr_346(8));
E(164)<=not ( sumr_347(0) or sumr_347(1) or sumr_347(2) or sumr_347(3) or sumr_347(4) or sumr_347(5) or sumr_347(6) or sumr_347(7) or sumr_347(8));
E(163)<=not ( sumr_348(0) or sumr_348(1) or sumr_348(2) or sumr_348(3) or sumr_348(4) or sumr_348(5) or sumr_348(6) or sumr_348(7) or sumr_348(8));
E(162)<=not ( sumr_349(0) or sumr_349(1) or sumr_349(2) or sumr_349(3) or sumr_349(4) or sumr_349(5) or sumr_349(6) or sumr_349(7) or sumr_349(8));
E(161)<=not ( sumr_350(0) or sumr_350(1) or sumr_350(2) or sumr_350(3) or sumr_350(4) or sumr_350(5) or sumr_350(6) or sumr_350(7) or sumr_350(8));
E(160)<=not ( sumr_351(0) or sumr_351(1) or sumr_351(2) or sumr_351(3) or sumr_351(4) or sumr_351(5) or sumr_351(6) or sumr_351(7) or sumr_351(8));
E(159)<=not ( sumr_352(0) or sumr_352(1) or sumr_352(2) or sumr_352(3) or sumr_352(4) or sumr_352(5) or sumr_352(6) or sumr_352(7) or sumr_352(8));
E(158)<=not ( sumr_353(0) or sumr_353(1) or sumr_353(2) or sumr_353(3) or sumr_353(4) or sumr_353(5) or sumr_353(6) or sumr_353(7) or sumr_353(8));
E(157)<=not ( sumr_354(0) or sumr_354(1) or sumr_354(2) or sumr_354(3) or sumr_354(4) or sumr_354(5) or sumr_354(6) or sumr_354(7) or sumr_354(8));
E(156)<=not ( sumr_355(0) or sumr_355(1) or sumr_355(2) or sumr_355(3) or sumr_355(4) or sumr_355(5) or sumr_355(6) or sumr_355(7) or sumr_355(8));
E(155)<=not ( sumr_356(0) or sumr_356(1) or sumr_356(2) or sumr_356(3) or sumr_356(4) or sumr_356(5) or sumr_356(6) or sumr_356(7) or sumr_356(8));
E(154)<=not ( sumr_357(0) or sumr_357(1) or sumr_357(2) or sumr_357(3) or sumr_357(4) or sumr_357(5) or sumr_357(6) or sumr_357(7) or sumr_357(8));
E(153)<=not ( sumr_358(0) or sumr_358(1) or sumr_358(2) or sumr_358(3) or sumr_358(4) or sumr_358(5) or sumr_358(6) or sumr_358(7) or sumr_358(8));
E(152)<=not ( sumr_359(0) or sumr_359(1) or sumr_359(2) or sumr_359(3) or sumr_359(4) or sumr_359(5) or sumr_359(6) or sumr_359(7) or sumr_359(8));
E(151)<=not ( sumr_360(0) or sumr_360(1) or sumr_360(2) or sumr_360(3) or sumr_360(4) or sumr_360(5) or sumr_360(6) or sumr_360(7) or sumr_360(8));
E(150)<=not ( sumr_361(0) or sumr_361(1) or sumr_361(2) or sumr_361(3) or sumr_361(4) or sumr_361(5) or sumr_361(6) or sumr_361(7) or sumr_361(8));
E(149)<=not ( sumr_362(0) or sumr_362(1) or sumr_362(2) or sumr_362(3) or sumr_362(4) or sumr_362(5) or sumr_362(6) or sumr_362(7) or sumr_362(8));
E(148)<=not ( sumr_363(0) or sumr_363(1) or sumr_363(2) or sumr_363(3) or sumr_363(4) or sumr_363(5) or sumr_363(6) or sumr_363(7) or sumr_363(8));
E(147)<=not ( sumr_364(0) or sumr_364(1) or sumr_364(2) or sumr_364(3) or sumr_364(4) or sumr_364(5) or sumr_364(6) or sumr_364(7) or sumr_364(8));
E(146)<=not ( sumr_365(0) or sumr_365(1) or sumr_365(2) or sumr_365(3) or sumr_365(4) or sumr_365(5) or sumr_365(6) or sumr_365(7) or sumr_365(8));
E(145)<=not ( sumr_366(0) or sumr_366(1) or sumr_366(2) or sumr_366(3) or sumr_366(4) or sumr_366(5) or sumr_366(6) or sumr_366(7) or sumr_366(8));
E(144)<=not ( sumr_367(0) or sumr_367(1) or sumr_367(2) or sumr_367(3) or sumr_367(4) or sumr_367(5) or sumr_367(6) or sumr_367(7) or sumr_367(8));
E(143)<=not ( sumr_368(0) or sumr_368(1) or sumr_368(2) or sumr_368(3) or sumr_368(4) or sumr_368(5) or sumr_368(6) or sumr_368(7) or sumr_368(8));
E(142)<=not ( sumr_369(0) or sumr_369(1) or sumr_369(2) or sumr_369(3) or sumr_369(4) or sumr_369(5) or sumr_369(6) or sumr_369(7) or sumr_369(8));
E(141)<=not ( sumr_370(0) or sumr_370(1) or sumr_370(2) or sumr_370(3) or sumr_370(4) or sumr_370(5) or sumr_370(6) or sumr_370(7) or sumr_370(8));
E(140)<=not ( sumr_371(0) or sumr_371(1) or sumr_371(2) or sumr_371(3) or sumr_371(4) or sumr_371(5) or sumr_371(6) or sumr_371(7) or sumr_371(8));
E(139)<=not ( sumr_372(0) or sumr_372(1) or sumr_372(2) or sumr_372(3) or sumr_372(4) or sumr_372(5) or sumr_372(6) or sumr_372(7) or sumr_372(8));
E(138)<=not ( sumr_373(0) or sumr_373(1) or sumr_373(2) or sumr_373(3) or sumr_373(4) or sumr_373(5) or sumr_373(6) or sumr_373(7) or sumr_373(8));
E(137)<=not ( sumr_374(0) or sumr_374(1) or sumr_374(2) or sumr_374(3) or sumr_374(4) or sumr_374(5) or sumr_374(6) or sumr_374(7) or sumr_374(8));
E(136)<=not ( sumr_375(0) or sumr_375(1) or sumr_375(2) or sumr_375(3) or sumr_375(4) or sumr_375(5) or sumr_375(6) or sumr_375(7) or sumr_375(8));
E(135)<=not ( sumr_376(0) or sumr_376(1) or sumr_376(2) or sumr_376(3) or sumr_376(4) or sumr_376(5) or sumr_376(6) or sumr_376(7) or sumr_376(8));
E(134)<=not ( sumr_377(0) or sumr_377(1) or sumr_377(2) or sumr_377(3) or sumr_377(4) or sumr_377(5) or sumr_377(6) or sumr_377(7) or sumr_377(8));
E(133)<=not ( sumr_378(0) or sumr_378(1) or sumr_378(2) or sumr_378(3) or sumr_378(4) or sumr_378(5) or sumr_378(6) or sumr_378(7) or sumr_378(8));
E(132)<=not ( sumr_379(0) or sumr_379(1) or sumr_379(2) or sumr_379(3) or sumr_379(4) or sumr_379(5) or sumr_379(6) or sumr_379(7) or sumr_379(8));
E(131)<=not ( sumr_380(0) or sumr_380(1) or sumr_380(2) or sumr_380(3) or sumr_380(4) or sumr_380(5) or sumr_380(6) or sumr_380(7) or sumr_380(8));
E(130)<=not ( sumr_381(0) or sumr_381(1) or sumr_381(2) or sumr_381(3) or sumr_381(4) or sumr_381(5) or sumr_381(6) or sumr_381(7) or sumr_381(8));
E(129)<=not ( sumr_382(0) or sumr_382(1) or sumr_382(2) or sumr_382(3) or sumr_382(4) or sumr_382(5) or sumr_382(6) or sumr_382(7) or sumr_382(8));
E(128)<=not ( sumr_383(0) or sumr_383(1) or sumr_383(2) or sumr_383(3) or sumr_383(4) or sumr_383(5) or sumr_383(6) or sumr_383(7) or sumr_383(8));
E(127)<=not ( sumr_384(0) or sumr_384(1) or sumr_384(2) or sumr_384(3) or sumr_384(4) or sumr_384(5) or sumr_384(6) or sumr_384(7) or sumr_384(8));
E(126)<=not ( sumr_385(0) or sumr_385(1) or sumr_385(2) or sumr_385(3) or sumr_385(4) or sumr_385(5) or sumr_385(6) or sumr_385(7) or sumr_385(8));
E(125)<=not ( sumr_386(0) or sumr_386(1) or sumr_386(2) or sumr_386(3) or sumr_386(4) or sumr_386(5) or sumr_386(6) or sumr_386(7) or sumr_386(8));
E(124)<=not ( sumr_387(0) or sumr_387(1) or sumr_387(2) or sumr_387(3) or sumr_387(4) or sumr_387(5) or sumr_387(6) or sumr_387(7) or sumr_387(8));
E(123)<=not ( sumr_388(0) or sumr_388(1) or sumr_388(2) or sumr_388(3) or sumr_388(4) or sumr_388(5) or sumr_388(6) or sumr_388(7) or sumr_388(8));
E(122)<=not ( sumr_389(0) or sumr_389(1) or sumr_389(2) or sumr_389(3) or sumr_389(4) or sumr_389(5) or sumr_389(6) or sumr_389(7) or sumr_389(8));
E(121)<=not ( sumr_390(0) or sumr_390(1) or sumr_390(2) or sumr_390(3) or sumr_390(4) or sumr_390(5) or sumr_390(6) or sumr_390(7) or sumr_390(8));
E(120)<=not ( sumr_391(0) or sumr_391(1) or sumr_391(2) or sumr_391(3) or sumr_391(4) or sumr_391(5) or sumr_391(6) or sumr_391(7) or sumr_391(8));
E(119)<=not ( sumr_392(0) or sumr_392(1) or sumr_392(2) or sumr_392(3) or sumr_392(4) or sumr_392(5) or sumr_392(6) or sumr_392(7) or sumr_392(8));
E(118)<=not ( sumr_393(0) or sumr_393(1) or sumr_393(2) or sumr_393(3) or sumr_393(4) or sumr_393(5) or sumr_393(6) or sumr_393(7) or sumr_393(8));
E(117)<=not ( sumr_394(0) or sumr_394(1) or sumr_394(2) or sumr_394(3) or sumr_394(4) or sumr_394(5) or sumr_394(6) or sumr_394(7) or sumr_394(8));
E(116)<=not ( sumr_395(0) or sumr_395(1) or sumr_395(2) or sumr_395(3) or sumr_395(4) or sumr_395(5) or sumr_395(6) or sumr_395(7) or sumr_395(8));
E(115)<=not ( sumr_396(0) or sumr_396(1) or sumr_396(2) or sumr_396(3) or sumr_396(4) or sumr_396(5) or sumr_396(6) or sumr_396(7) or sumr_396(8));
E(114)<=not ( sumr_397(0) or sumr_397(1) or sumr_397(2) or sumr_397(3) or sumr_397(4) or sumr_397(5) or sumr_397(6) or sumr_397(7) or sumr_397(8));
E(113)<=not ( sumr_398(0) or sumr_398(1) or sumr_398(2) or sumr_398(3) or sumr_398(4) or sumr_398(5) or sumr_398(6) or sumr_398(7) or sumr_398(8));
E(112)<=not ( sumr_399(0) or sumr_399(1) or sumr_399(2) or sumr_399(3) or sumr_399(4) or sumr_399(5) or sumr_399(6) or sumr_399(7) or sumr_399(8));
E(111)<=not ( sumr_400(0) or sumr_400(1) or sumr_400(2) or sumr_400(3) or sumr_400(4) or sumr_400(5) or sumr_400(6) or sumr_400(7) or sumr_400(8));
E(110)<=not ( sumr_401(0) or sumr_401(1) or sumr_401(2) or sumr_401(3) or sumr_401(4) or sumr_401(5) or sumr_401(6) or sumr_401(7) or sumr_401(8));
E(109)<=not ( sumr_402(0) or sumr_402(1) or sumr_402(2) or sumr_402(3) or sumr_402(4) or sumr_402(5) or sumr_402(6) or sumr_402(7) or sumr_402(8));
E(108)<=not ( sumr_403(0) or sumr_403(1) or sumr_403(2) or sumr_403(3) or sumr_403(4) or sumr_403(5) or sumr_403(6) or sumr_403(7) or sumr_403(8));
E(107)<=not ( sumr_404(0) or sumr_404(1) or sumr_404(2) or sumr_404(3) or sumr_404(4) or sumr_404(5) or sumr_404(6) or sumr_404(7) or sumr_404(8));
E(106)<=not ( sumr_405(0) or sumr_405(1) or sumr_405(2) or sumr_405(3) or sumr_405(4) or sumr_405(5) or sumr_405(6) or sumr_405(7) or sumr_405(8));
E(105)<=not ( sumr_406(0) or sumr_406(1) or sumr_406(2) or sumr_406(3) or sumr_406(4) or sumr_406(5) or sumr_406(6) or sumr_406(7) or sumr_406(8));
E(104)<=not ( sumr_407(0) or sumr_407(1) or sumr_407(2) or sumr_407(3) or sumr_407(4) or sumr_407(5) or sumr_407(6) or sumr_407(7) or sumr_407(8));
E(103)<=not ( sumr_408(0) or sumr_408(1) or sumr_408(2) or sumr_408(3) or sumr_408(4) or sumr_408(5) or sumr_408(6) or sumr_408(7) or sumr_408(8));
E(102)<=not ( sumr_409(0) or sumr_409(1) or sumr_409(2) or sumr_409(3) or sumr_409(4) or sumr_409(5) or sumr_409(6) or sumr_409(7) or sumr_409(8));
E(101)<=not ( sumr_410(0) or sumr_410(1) or sumr_410(2) or sumr_410(3) or sumr_410(4) or sumr_410(5) or sumr_410(6) or sumr_410(7) or sumr_410(8));
E(100)<=not ( sumr_411(0) or sumr_411(1) or sumr_411(2) or sumr_411(3) or sumr_411(4) or sumr_411(5) or sumr_411(6) or sumr_411(7) or sumr_411(8));
E(99)<=not ( sumr_412(0) or sumr_412(1) or sumr_412(2) or sumr_412(3) or sumr_412(4) or sumr_412(5) or sumr_412(6) or sumr_412(7) or sumr_412(8));
E(98)<=not ( sumr_413(0) or sumr_413(1) or sumr_413(2) or sumr_413(3) or sumr_413(4) or sumr_413(5) or sumr_413(6) or sumr_413(7) or sumr_413(8));
E(97)<=not ( sumr_414(0) or sumr_414(1) or sumr_414(2) or sumr_414(3) or sumr_414(4) or sumr_414(5) or sumr_414(6) or sumr_414(7) or sumr_414(8));
E(96)<=not ( sumr_415(0) or sumr_415(1) or sumr_415(2) or sumr_415(3) or sumr_415(4) or sumr_415(5) or sumr_415(6) or sumr_415(7) or sumr_415(8));
E(95)<=not ( sumr_416(0) or sumr_416(1) or sumr_416(2) or sumr_416(3) or sumr_416(4) or sumr_416(5) or sumr_416(6) or sumr_416(7) or sumr_416(8));
E(94)<=not ( sumr_417(0) or sumr_417(1) or sumr_417(2) or sumr_417(3) or sumr_417(4) or sumr_417(5) or sumr_417(6) or sumr_417(7) or sumr_417(8));
E(93)<=not ( sumr_418(0) or sumr_418(1) or sumr_418(2) or sumr_418(3) or sumr_418(4) or sumr_418(5) or sumr_418(6) or sumr_418(7) or sumr_418(8));
E(92)<=not ( sumr_419(0) or sumr_419(1) or sumr_419(2) or sumr_419(3) or sumr_419(4) or sumr_419(5) or sumr_419(6) or sumr_419(7) or sumr_419(8));
E(91)<=not ( sumr_420(0) or sumr_420(1) or sumr_420(2) or sumr_420(3) or sumr_420(4) or sumr_420(5) or sumr_420(6) or sumr_420(7) or sumr_420(8));
E(90)<=not ( sumr_421(0) or sumr_421(1) or sumr_421(2) or sumr_421(3) or sumr_421(4) or sumr_421(5) or sumr_421(6) or sumr_421(7) or sumr_421(8));
E(89)<=not ( sumr_422(0) or sumr_422(1) or sumr_422(2) or sumr_422(3) or sumr_422(4) or sumr_422(5) or sumr_422(6) or sumr_422(7) or sumr_422(8));
E(88)<=not ( sumr_423(0) or sumr_423(1) or sumr_423(2) or sumr_423(3) or sumr_423(4) or sumr_423(5) or sumr_423(6) or sumr_423(7) or sumr_423(8));
E(87)<=not ( sumr_424(0) or sumr_424(1) or sumr_424(2) or sumr_424(3) or sumr_424(4) or sumr_424(5) or sumr_424(6) or sumr_424(7) or sumr_424(8));
E(86)<=not ( sumr_425(0) or sumr_425(1) or sumr_425(2) or sumr_425(3) or sumr_425(4) or sumr_425(5) or sumr_425(6) or sumr_425(7) or sumr_425(8));
E(85)<=not ( sumr_426(0) or sumr_426(1) or sumr_426(2) or sumr_426(3) or sumr_426(4) or sumr_426(5) or sumr_426(6) or sumr_426(7) or sumr_426(8));
E(84)<=not ( sumr_427(0) or sumr_427(1) or sumr_427(2) or sumr_427(3) or sumr_427(4) or sumr_427(5) or sumr_427(6) or sumr_427(7) or sumr_427(8));
E(83)<=not ( sumr_428(0) or sumr_428(1) or sumr_428(2) or sumr_428(3) or sumr_428(4) or sumr_428(5) or sumr_428(6) or sumr_428(7) or sumr_428(8));
E(82)<=not ( sumr_429(0) or sumr_429(1) or sumr_429(2) or sumr_429(3) or sumr_429(4) or sumr_429(5) or sumr_429(6) or sumr_429(7) or sumr_429(8));
E(81)<=not ( sumr_430(0) or sumr_430(1) or sumr_430(2) or sumr_430(3) or sumr_430(4) or sumr_430(5) or sumr_430(6) or sumr_430(7) or sumr_430(8));
E(80)<=not ( sumr_431(0) or sumr_431(1) or sumr_431(2) or sumr_431(3) or sumr_431(4) or sumr_431(5) or sumr_431(6) or sumr_431(7) or sumr_431(8));
E(79)<=not ( sumr_432(0) or sumr_432(1) or sumr_432(2) or sumr_432(3) or sumr_432(4) or sumr_432(5) or sumr_432(6) or sumr_432(7) or sumr_432(8));
E(78)<=not ( sumr_433(0) or sumr_433(1) or sumr_433(2) or sumr_433(3) or sumr_433(4) or sumr_433(5) or sumr_433(6) or sumr_433(7) or sumr_433(8));
E(77)<=not ( sumr_434(0) or sumr_434(1) or sumr_434(2) or sumr_434(3) or sumr_434(4) or sumr_434(5) or sumr_434(6) or sumr_434(7) or sumr_434(8));
E(76)<=not ( sumr_435(0) or sumr_435(1) or sumr_435(2) or sumr_435(3) or sumr_435(4) or sumr_435(5) or sumr_435(6) or sumr_435(7) or sumr_435(8));
E(75)<=not ( sumr_436(0) or sumr_436(1) or sumr_436(2) or sumr_436(3) or sumr_436(4) or sumr_436(5) or sumr_436(6) or sumr_436(7) or sumr_436(8));
E(74)<=not ( sumr_437(0) or sumr_437(1) or sumr_437(2) or sumr_437(3) or sumr_437(4) or sumr_437(5) or sumr_437(6) or sumr_437(7) or sumr_437(8));
E(73)<=not ( sumr_438(0) or sumr_438(1) or sumr_438(2) or sumr_438(3) or sumr_438(4) or sumr_438(5) or sumr_438(6) or sumr_438(7) or sumr_438(8));
E(72)<=not ( sumr_439(0) or sumr_439(1) or sumr_439(2) or sumr_439(3) or sumr_439(4) or sumr_439(5) or sumr_439(6) or sumr_439(7) or sumr_439(8));
E(71)<=not ( sumr_440(0) or sumr_440(1) or sumr_440(2) or sumr_440(3) or sumr_440(4) or sumr_440(5) or sumr_440(6) or sumr_440(7) or sumr_440(8));
E(70)<=not ( sumr_441(0) or sumr_441(1) or sumr_441(2) or sumr_441(3) or sumr_441(4) or sumr_441(5) or sumr_441(6) or sumr_441(7) or sumr_441(8));
E(69)<=not ( sumr_442(0) or sumr_442(1) or sumr_442(2) or sumr_442(3) or sumr_442(4) or sumr_442(5) or sumr_442(6) or sumr_442(7) or sumr_442(8));
E(68)<=not ( sumr_443(0) or sumr_443(1) or sumr_443(2) or sumr_443(3) or sumr_443(4) or sumr_443(5) or sumr_443(6) or sumr_443(7) or sumr_443(8));
E(67)<=not ( sumr_444(0) or sumr_444(1) or sumr_444(2) or sumr_444(3) or sumr_444(4) or sumr_444(5) or sumr_444(6) or sumr_444(7) or sumr_444(8));
E(66)<=not ( sumr_445(0) or sumr_445(1) or sumr_445(2) or sumr_445(3) or sumr_445(4) or sumr_445(5) or sumr_445(6) or sumr_445(7) or sumr_445(8));
E(65)<=not ( sumr_446(0) or sumr_446(1) or sumr_446(2) or sumr_446(3) or sumr_446(4) or sumr_446(5) or sumr_446(6) or sumr_446(7) or sumr_446(8));
E(64)<=not ( sumr_447(0) or sumr_447(1) or sumr_447(2) or sumr_447(3) or sumr_447(4) or sumr_447(5) or sumr_447(6) or sumr_447(7) or sumr_447(8));
E(63)<=not ( sumr_448(0) or sumr_448(1) or sumr_448(2) or sumr_448(3) or sumr_448(4) or sumr_448(5) or sumr_448(6) or sumr_448(7) or sumr_448(8));
E(62)<=not ( sumr_449(0) or sumr_449(1) or sumr_449(2) or sumr_449(3) or sumr_449(4) or sumr_449(5) or sumr_449(6) or sumr_449(7) or sumr_449(8));
E(61)<=not ( sumr_450(0) or sumr_450(1) or sumr_450(2) or sumr_450(3) or sumr_450(4) or sumr_450(5) or sumr_450(6) or sumr_450(7) or sumr_450(8));
E(60)<=not ( sumr_451(0) or sumr_451(1) or sumr_451(2) or sumr_451(3) or sumr_451(4) or sumr_451(5) or sumr_451(6) or sumr_451(7) or sumr_451(8));
E(59)<=not ( sumr_452(0) or sumr_452(1) or sumr_452(2) or sumr_452(3) or sumr_452(4) or sumr_452(5) or sumr_452(6) or sumr_452(7) or sumr_452(8));
E(58)<=not ( sumr_453(0) or sumr_453(1) or sumr_453(2) or sumr_453(3) or sumr_453(4) or sumr_453(5) or sumr_453(6) or sumr_453(7) or sumr_453(8));
E(57)<=not ( sumr_454(0) or sumr_454(1) or sumr_454(2) or sumr_454(3) or sumr_454(4) or sumr_454(5) or sumr_454(6) or sumr_454(7) or sumr_454(8));
E(56)<=not ( sumr_455(0) or sumr_455(1) or sumr_455(2) or sumr_455(3) or sumr_455(4) or sumr_455(5) or sumr_455(6) or sumr_455(7) or sumr_455(8));
E(55)<=not ( sumr_456(0) or sumr_456(1) or sumr_456(2) or sumr_456(3) or sumr_456(4) or sumr_456(5) or sumr_456(6) or sumr_456(7) or sumr_456(8));
E(54)<=not ( sumr_457(0) or sumr_457(1) or sumr_457(2) or sumr_457(3) or sumr_457(4) or sumr_457(5) or sumr_457(6) or sumr_457(7) or sumr_457(8));
E(53)<=not ( sumr_458(0) or sumr_458(1) or sumr_458(2) or sumr_458(3) or sumr_458(4) or sumr_458(5) or sumr_458(6) or sumr_458(7) or sumr_458(8));
E(52)<=not ( sumr_459(0) or sumr_459(1) or sumr_459(2) or sumr_459(3) or sumr_459(4) or sumr_459(5) or sumr_459(6) or sumr_459(7) or sumr_459(8));
E(51)<=not ( sumr_460(0) or sumr_460(1) or sumr_460(2) or sumr_460(3) or sumr_460(4) or sumr_460(5) or sumr_460(6) or sumr_460(7) or sumr_460(8));
E(50)<=not ( sumr_461(0) or sumr_461(1) or sumr_461(2) or sumr_461(3) or sumr_461(4) or sumr_461(5) or sumr_461(6) or sumr_461(7) or sumr_461(8));
E(49)<=not ( sumr_462(0) or sumr_462(1) or sumr_462(2) or sumr_462(3) or sumr_462(4) or sumr_462(5) or sumr_462(6) or sumr_462(7) or sumr_462(8));
E(48)<=not ( sumr_463(0) or sumr_463(1) or sumr_463(2) or sumr_463(3) or sumr_463(4) or sumr_463(5) or sumr_463(6) or sumr_463(7) or sumr_463(8));
E(47)<=not ( sumr_464(0) or sumr_464(1) or sumr_464(2) or sumr_464(3) or sumr_464(4) or sumr_464(5) or sumr_464(6) or sumr_464(7) or sumr_464(8));
E(46)<=not ( sumr_465(0) or sumr_465(1) or sumr_465(2) or sumr_465(3) or sumr_465(4) or sumr_465(5) or sumr_465(6) or sumr_465(7) or sumr_465(8));
E(45)<=not ( sumr_466(0) or sumr_466(1) or sumr_466(2) or sumr_466(3) or sumr_466(4) or sumr_466(5) or sumr_466(6) or sumr_466(7) or sumr_466(8));
E(44)<=not ( sumr_467(0) or sumr_467(1) or sumr_467(2) or sumr_467(3) or sumr_467(4) or sumr_467(5) or sumr_467(6) or sumr_467(7) or sumr_467(8));
E(43)<=not ( sumr_468(0) or sumr_468(1) or sumr_468(2) or sumr_468(3) or sumr_468(4) or sumr_468(5) or sumr_468(6) or sumr_468(7) or sumr_468(8));
E(42)<=not ( sumr_469(0) or sumr_469(1) or sumr_469(2) or sumr_469(3) or sumr_469(4) or sumr_469(5) or sumr_469(6) or sumr_469(7) or sumr_469(8));
E(41)<=not ( sumr_470(0) or sumr_470(1) or sumr_470(2) or sumr_470(3) or sumr_470(4) or sumr_470(5) or sumr_470(6) or sumr_470(7) or sumr_470(8));
E(40)<=not ( sumr_471(0) or sumr_471(1) or sumr_471(2) or sumr_471(3) or sumr_471(4) or sumr_471(5) or sumr_471(6) or sumr_471(7) or sumr_471(8));
E(39)<=not ( sumr_472(0) or sumr_472(1) or sumr_472(2) or sumr_472(3) or sumr_472(4) or sumr_472(5) or sumr_472(6) or sumr_472(7) or sumr_472(8));
E(38)<=not ( sumr_473(0) or sumr_473(1) or sumr_473(2) or sumr_473(3) or sumr_473(4) or sumr_473(5) or sumr_473(6) or sumr_473(7) or sumr_473(8));
E(37)<=not ( sumr_474(0) or sumr_474(1) or sumr_474(2) or sumr_474(3) or sumr_474(4) or sumr_474(5) or sumr_474(6) or sumr_474(7) or sumr_474(8));
E(36)<=not ( sumr_475(0) or sumr_475(1) or sumr_475(2) or sumr_475(3) or sumr_475(4) or sumr_475(5) or sumr_475(6) or sumr_475(7) or sumr_475(8));
E(35)<=not ( sumr_476(0) or sumr_476(1) or sumr_476(2) or sumr_476(3) or sumr_476(4) or sumr_476(5) or sumr_476(6) or sumr_476(7) or sumr_476(8));
E(34)<=not ( sumr_477(0) or sumr_477(1) or sumr_477(2) or sumr_477(3) or sumr_477(4) or sumr_477(5) or sumr_477(6) or sumr_477(7) or sumr_477(8));
E(33)<=not ( sumr_478(0) or sumr_478(1) or sumr_478(2) or sumr_478(3) or sumr_478(4) or sumr_478(5) or sumr_478(6) or sumr_478(7) or sumr_478(8));
E(32)<=not ( sumr_479(0) or sumr_479(1) or sumr_479(2) or sumr_479(3) or sumr_479(4) or sumr_479(5) or sumr_479(6) or sumr_479(7) or sumr_479(8));
E(31)<=not ( sumr_480(0) or sumr_480(1) or sumr_480(2) or sumr_480(3) or sumr_480(4) or sumr_480(5) or sumr_480(6) or sumr_480(7) or sumr_480(8));
E(30)<=not ( sumr_481(0) or sumr_481(1) or sumr_481(2) or sumr_481(3) or sumr_481(4) or sumr_481(5) or sumr_481(6) or sumr_481(7) or sumr_481(8));
E(29)<=not ( sumr_482(0) or sumr_482(1) or sumr_482(2) or sumr_482(3) or sumr_482(4) or sumr_482(5) or sumr_482(6) or sumr_482(7) or sumr_482(8));
E(28)<=not ( sumr_483(0) or sumr_483(1) or sumr_483(2) or sumr_483(3) or sumr_483(4) or sumr_483(5) or sumr_483(6) or sumr_483(7) or sumr_483(8));
E(27)<=not ( sumr_484(0) or sumr_484(1) or sumr_484(2) or sumr_484(3) or sumr_484(4) or sumr_484(5) or sumr_484(6) or sumr_484(7) or sumr_484(8));
E(26)<=not ( sumr_485(0) or sumr_485(1) or sumr_485(2) or sumr_485(3) or sumr_485(4) or sumr_485(5) or sumr_485(6) or sumr_485(7) or sumr_485(8));
E(25)<=not ( sumr_486(0) or sumr_486(1) or sumr_486(2) or sumr_486(3) or sumr_486(4) or sumr_486(5) or sumr_486(6) or sumr_486(7) or sumr_486(8));
E(24)<=not ( sumr_487(0) or sumr_487(1) or sumr_487(2) or sumr_487(3) or sumr_487(4) or sumr_487(5) or sumr_487(6) or sumr_487(7) or sumr_487(8));
E(23)<=not ( sumr_488(0) or sumr_488(1) or sumr_488(2) or sumr_488(3) or sumr_488(4) or sumr_488(5) or sumr_488(6) or sumr_488(7) or sumr_488(8));
E(22)<=not ( sumr_489(0) or sumr_489(1) or sumr_489(2) or sumr_489(3) or sumr_489(4) or sumr_489(5) or sumr_489(6) or sumr_489(7) or sumr_489(8));
E(21)<=not ( sumr_490(0) or sumr_490(1) or sumr_490(2) or sumr_490(3) or sumr_490(4) or sumr_490(5) or sumr_490(6) or sumr_490(7) or sumr_490(8));
E(20)<=not ( sumr_491(0) or sumr_491(1) or sumr_491(2) or sumr_491(3) or sumr_491(4) or sumr_491(5) or sumr_491(6) or sumr_491(7) or sumr_491(8));
E(19)<=not ( sumr_492(0) or sumr_492(1) or sumr_492(2) or sumr_492(3) or sumr_492(4) or sumr_492(5) or sumr_492(6) or sumr_492(7) or sumr_492(8));
E(18)<=not ( sumr_493(0) or sumr_493(1) or sumr_493(2) or sumr_493(3) or sumr_493(4) or sumr_493(5) or sumr_493(6) or sumr_493(7) or sumr_493(8));
E(17)<=not ( sumr_494(0) or sumr_494(1) or sumr_494(2) or sumr_494(3) or sumr_494(4) or sumr_494(5) or sumr_494(6) or sumr_494(7) or sumr_494(8));
E(16)<=not ( sumr_495(0) or sumr_495(1) or sumr_495(2) or sumr_495(3) or sumr_495(4) or sumr_495(5) or sumr_495(6) or sumr_495(7) or sumr_495(8));
E(15)<=not ( sumr_496(0) or sumr_496(1) or sumr_496(2) or sumr_496(3) or sumr_496(4) or sumr_496(5) or sumr_496(6) or sumr_496(7) or sumr_496(8));
E(14)<=not ( sumr_497(0) or sumr_497(1) or sumr_497(2) or sumr_497(3) or sumr_497(4) or sumr_497(5) or sumr_497(6) or sumr_497(7) or sumr_497(8));
E(13)<=not ( sumr_498(0) or sumr_498(1) or sumr_498(2) or sumr_498(3) or sumr_498(4) or sumr_498(5) or sumr_498(6) or sumr_498(7) or sumr_498(8));
E(12)<=not ( sumr_499(0) or sumr_499(1) or sumr_499(2) or sumr_499(3) or sumr_499(4) or sumr_499(5) or sumr_499(6) or sumr_499(7) or sumr_499(8));
E(11)<=not ( sumr_500(0) or sumr_500(1) or sumr_500(2) or sumr_500(3) or sumr_500(4) or sumr_500(5) or sumr_500(6) or sumr_500(7) or sumr_500(8));
E(10)<=not ( sumr_501(0) or sumr_501(1) or sumr_501(2) or sumr_501(3) or sumr_501(4) or sumr_501(5) or sumr_501(6) or sumr_501(7) or sumr_501(8));
E(9)<=not ( sumr_502(0) or sumr_502(1) or sumr_502(2) or sumr_502(3) or sumr_502(4) or sumr_502(5) or sumr_502(6) or sumr_502(7) or sumr_502(8));
E(8)<=not ( sumr_503(0) or sumr_503(1) or sumr_503(2) or sumr_503(3) or sumr_503(4) or sumr_503(5) or sumr_503(6) or sumr_503(7) or sumr_503(8));
E(7)<=not ( sumr_504(0) or sumr_504(1) or sumr_504(2) or sumr_504(3) or sumr_504(4) or sumr_504(5) or sumr_504(6) or sumr_504(7) or sumr_504(8));
E(6)<=not ( sumr_505(0) or sumr_505(1) or sumr_505(2) or sumr_505(3) or sumr_505(4) or sumr_505(5) or sumr_505(6) or sumr_505(7) or sumr_505(8));
E(5)<=not ( sumr_506(0) or sumr_506(1) or sumr_506(2) or sumr_506(3) or sumr_506(4) or sumr_506(5) or sumr_506(6) or sumr_506(7) or sumr_506(8));
E(4)<=not ( sumr_507(0) or sumr_507(1) or sumr_507(2) or sumr_507(3) or sumr_507(4) or sumr_507(5) or sumr_507(6) or sumr_507(7) or sumr_507(8));
E(3)<=not ( sumr_508(0) or sumr_508(1) or sumr_508(2) or sumr_508(3) or sumr_508(4) or sumr_508(5) or sumr_508(6) or sumr_508(7) or sumr_508(8));
E(2)<=not ( sumr_509(0) or sumr_509(1) or sumr_509(2) or sumr_509(3) or sumr_509(4) or sumr_509(5) or sumr_509(6) or sumr_509(7) or sumr_509(8));
E(1)<=not ( sumr_510(0) or sumr_510(1) or sumr_510(2) or sumr_510(3) or sumr_510(4) or sumr_510(5) or sumr_510(6) or sumr_510(7) or sumr_510(8));
E(0)<=not ( sumr_511(0) or sumr_511(1) or sumr_511(2) or sumr_511(3) or sumr_511(4) or sumr_511(5) or sumr_511(6) or sumr_511(7) or sumr_511(8));
end arch;
