library ieee;
use ieee.std_logic_1164.all;
entity chien is
    port(
        a_1     :    in  std_logic_vector(7 downto 0);
        a_2     :    in  std_logic_vector(7 downto 0);
        E     :    out std_logic_vector(254 downto 0)
);
end entity;

architecture arch of chien is
    signal mulr_1_1 : std_logic_vector(7 downto 0);
    signal mulr_2_1 : std_logic_vector(7 downto 0);
    signal mulr_1_2 : std_logic_vector(7 downto 0);
    signal mulr_2_2 : std_logic_vector(7 downto 0);
    signal mulr_1_3 : std_logic_vector(7 downto 0);
    signal mulr_2_3 : std_logic_vector(7 downto 0);
    signal mulr_1_4 : std_logic_vector(7 downto 0);
    signal mulr_2_4 : std_logic_vector(7 downto 0);
    signal mulr_1_5 : std_logic_vector(7 downto 0);
    signal mulr_2_5 : std_logic_vector(7 downto 0);
    signal mulr_1_6 : std_logic_vector(7 downto 0);
    signal mulr_2_6 : std_logic_vector(7 downto 0);
    signal mulr_1_7 : std_logic_vector(7 downto 0);
    signal mulr_2_7 : std_logic_vector(7 downto 0);
    signal mulr_1_8 : std_logic_vector(7 downto 0);
    signal mulr_2_8 : std_logic_vector(7 downto 0);
    signal mulr_1_9 : std_logic_vector(7 downto 0);
    signal mulr_2_9 : std_logic_vector(7 downto 0);
    signal mulr_1_10 : std_logic_vector(7 downto 0);
    signal mulr_2_10 : std_logic_vector(7 downto 0);
    signal mulr_1_11 : std_logic_vector(7 downto 0);
    signal mulr_2_11 : std_logic_vector(7 downto 0);
    signal mulr_1_12 : std_logic_vector(7 downto 0);
    signal mulr_2_12 : std_logic_vector(7 downto 0);
    signal mulr_1_13 : std_logic_vector(7 downto 0);
    signal mulr_2_13 : std_logic_vector(7 downto 0);
    signal mulr_1_14 : std_logic_vector(7 downto 0);
    signal mulr_2_14 : std_logic_vector(7 downto 0);
    signal mulr_1_15 : std_logic_vector(7 downto 0);
    signal mulr_2_15 : std_logic_vector(7 downto 0);
    signal mulr_1_16 : std_logic_vector(7 downto 0);
    signal mulr_2_16 : std_logic_vector(7 downto 0);
    signal mulr_1_17 : std_logic_vector(7 downto 0);
    signal mulr_2_17 : std_logic_vector(7 downto 0);
    signal mulr_1_18 : std_logic_vector(7 downto 0);
    signal mulr_2_18 : std_logic_vector(7 downto 0);
    signal mulr_1_19 : std_logic_vector(7 downto 0);
    signal mulr_2_19 : std_logic_vector(7 downto 0);
    signal mulr_1_20 : std_logic_vector(7 downto 0);
    signal mulr_2_20 : std_logic_vector(7 downto 0);
    signal mulr_1_21 : std_logic_vector(7 downto 0);
    signal mulr_2_21 : std_logic_vector(7 downto 0);
    signal mulr_1_22 : std_logic_vector(7 downto 0);
    signal mulr_2_22 : std_logic_vector(7 downto 0);
    signal mulr_1_23 : std_logic_vector(7 downto 0);
    signal mulr_2_23 : std_logic_vector(7 downto 0);
    signal mulr_1_24 : std_logic_vector(7 downto 0);
    signal mulr_2_24 : std_logic_vector(7 downto 0);
    signal mulr_1_25 : std_logic_vector(7 downto 0);
    signal mulr_2_25 : std_logic_vector(7 downto 0);
    signal mulr_1_26 : std_logic_vector(7 downto 0);
    signal mulr_2_26 : std_logic_vector(7 downto 0);
    signal mulr_1_27 : std_logic_vector(7 downto 0);
    signal mulr_2_27 : std_logic_vector(7 downto 0);
    signal mulr_1_28 : std_logic_vector(7 downto 0);
    signal mulr_2_28 : std_logic_vector(7 downto 0);
    signal mulr_1_29 : std_logic_vector(7 downto 0);
    signal mulr_2_29 : std_logic_vector(7 downto 0);
    signal mulr_1_30 : std_logic_vector(7 downto 0);
    signal mulr_2_30 : std_logic_vector(7 downto 0);
    signal mulr_1_31 : std_logic_vector(7 downto 0);
    signal mulr_2_31 : std_logic_vector(7 downto 0);
    signal mulr_1_32 : std_logic_vector(7 downto 0);
    signal mulr_2_32 : std_logic_vector(7 downto 0);
    signal mulr_1_33 : std_logic_vector(7 downto 0);
    signal mulr_2_33 : std_logic_vector(7 downto 0);
    signal mulr_1_34 : std_logic_vector(7 downto 0);
    signal mulr_2_34 : std_logic_vector(7 downto 0);
    signal mulr_1_35 : std_logic_vector(7 downto 0);
    signal mulr_2_35 : std_logic_vector(7 downto 0);
    signal mulr_1_36 : std_logic_vector(7 downto 0);
    signal mulr_2_36 : std_logic_vector(7 downto 0);
    signal mulr_1_37 : std_logic_vector(7 downto 0);
    signal mulr_2_37 : std_logic_vector(7 downto 0);
    signal mulr_1_38 : std_logic_vector(7 downto 0);
    signal mulr_2_38 : std_logic_vector(7 downto 0);
    signal mulr_1_39 : std_logic_vector(7 downto 0);
    signal mulr_2_39 : std_logic_vector(7 downto 0);
    signal mulr_1_40 : std_logic_vector(7 downto 0);
    signal mulr_2_40 : std_logic_vector(7 downto 0);
    signal mulr_1_41 : std_logic_vector(7 downto 0);
    signal mulr_2_41 : std_logic_vector(7 downto 0);
    signal mulr_1_42 : std_logic_vector(7 downto 0);
    signal mulr_2_42 : std_logic_vector(7 downto 0);
    signal mulr_1_43 : std_logic_vector(7 downto 0);
    signal mulr_2_43 : std_logic_vector(7 downto 0);
    signal mulr_1_44 : std_logic_vector(7 downto 0);
    signal mulr_2_44 : std_logic_vector(7 downto 0);
    signal mulr_1_45 : std_logic_vector(7 downto 0);
    signal mulr_2_45 : std_logic_vector(7 downto 0);
    signal mulr_1_46 : std_logic_vector(7 downto 0);
    signal mulr_2_46 : std_logic_vector(7 downto 0);
    signal mulr_1_47 : std_logic_vector(7 downto 0);
    signal mulr_2_47 : std_logic_vector(7 downto 0);
    signal mulr_1_48 : std_logic_vector(7 downto 0);
    signal mulr_2_48 : std_logic_vector(7 downto 0);
    signal mulr_1_49 : std_logic_vector(7 downto 0);
    signal mulr_2_49 : std_logic_vector(7 downto 0);
    signal mulr_1_50 : std_logic_vector(7 downto 0);
    signal mulr_2_50 : std_logic_vector(7 downto 0);
    signal mulr_1_51 : std_logic_vector(7 downto 0);
    signal mulr_2_51 : std_logic_vector(7 downto 0);
    signal mulr_1_52 : std_logic_vector(7 downto 0);
    signal mulr_2_52 : std_logic_vector(7 downto 0);
    signal mulr_1_53 : std_logic_vector(7 downto 0);
    signal mulr_2_53 : std_logic_vector(7 downto 0);
    signal mulr_1_54 : std_logic_vector(7 downto 0);
    signal mulr_2_54 : std_logic_vector(7 downto 0);
    signal mulr_1_55 : std_logic_vector(7 downto 0);
    signal mulr_2_55 : std_logic_vector(7 downto 0);
    signal mulr_1_56 : std_logic_vector(7 downto 0);
    signal mulr_2_56 : std_logic_vector(7 downto 0);
    signal mulr_1_57 : std_logic_vector(7 downto 0);
    signal mulr_2_57 : std_logic_vector(7 downto 0);
    signal mulr_1_58 : std_logic_vector(7 downto 0);
    signal mulr_2_58 : std_logic_vector(7 downto 0);
    signal mulr_1_59 : std_logic_vector(7 downto 0);
    signal mulr_2_59 : std_logic_vector(7 downto 0);
    signal mulr_1_60 : std_logic_vector(7 downto 0);
    signal mulr_2_60 : std_logic_vector(7 downto 0);
    signal mulr_1_61 : std_logic_vector(7 downto 0);
    signal mulr_2_61 : std_logic_vector(7 downto 0);
    signal mulr_1_62 : std_logic_vector(7 downto 0);
    signal mulr_2_62 : std_logic_vector(7 downto 0);
    signal mulr_1_63 : std_logic_vector(7 downto 0);
    signal mulr_2_63 : std_logic_vector(7 downto 0);
    signal mulr_1_64 : std_logic_vector(7 downto 0);
    signal mulr_2_64 : std_logic_vector(7 downto 0);
    signal mulr_1_65 : std_logic_vector(7 downto 0);
    signal mulr_2_65 : std_logic_vector(7 downto 0);
    signal mulr_1_66 : std_logic_vector(7 downto 0);
    signal mulr_2_66 : std_logic_vector(7 downto 0);
    signal mulr_1_67 : std_logic_vector(7 downto 0);
    signal mulr_2_67 : std_logic_vector(7 downto 0);
    signal mulr_1_68 : std_logic_vector(7 downto 0);
    signal mulr_2_68 : std_logic_vector(7 downto 0);
    signal mulr_1_69 : std_logic_vector(7 downto 0);
    signal mulr_2_69 : std_logic_vector(7 downto 0);
    signal mulr_1_70 : std_logic_vector(7 downto 0);
    signal mulr_2_70 : std_logic_vector(7 downto 0);
    signal mulr_1_71 : std_logic_vector(7 downto 0);
    signal mulr_2_71 : std_logic_vector(7 downto 0);
    signal mulr_1_72 : std_logic_vector(7 downto 0);
    signal mulr_2_72 : std_logic_vector(7 downto 0);
    signal mulr_1_73 : std_logic_vector(7 downto 0);
    signal mulr_2_73 : std_logic_vector(7 downto 0);
    signal mulr_1_74 : std_logic_vector(7 downto 0);
    signal mulr_2_74 : std_logic_vector(7 downto 0);
    signal mulr_1_75 : std_logic_vector(7 downto 0);
    signal mulr_2_75 : std_logic_vector(7 downto 0);
    signal mulr_1_76 : std_logic_vector(7 downto 0);
    signal mulr_2_76 : std_logic_vector(7 downto 0);
    signal mulr_1_77 : std_logic_vector(7 downto 0);
    signal mulr_2_77 : std_logic_vector(7 downto 0);
    signal mulr_1_78 : std_logic_vector(7 downto 0);
    signal mulr_2_78 : std_logic_vector(7 downto 0);
    signal mulr_1_79 : std_logic_vector(7 downto 0);
    signal mulr_2_79 : std_logic_vector(7 downto 0);
    signal mulr_1_80 : std_logic_vector(7 downto 0);
    signal mulr_2_80 : std_logic_vector(7 downto 0);
    signal mulr_1_81 : std_logic_vector(7 downto 0);
    signal mulr_2_81 : std_logic_vector(7 downto 0);
    signal mulr_1_82 : std_logic_vector(7 downto 0);
    signal mulr_2_82 : std_logic_vector(7 downto 0);
    signal mulr_1_83 : std_logic_vector(7 downto 0);
    signal mulr_2_83 : std_logic_vector(7 downto 0);
    signal mulr_1_84 : std_logic_vector(7 downto 0);
    signal mulr_2_84 : std_logic_vector(7 downto 0);
    signal mulr_1_85 : std_logic_vector(7 downto 0);
    signal mulr_2_85 : std_logic_vector(7 downto 0);
    signal mulr_1_86 : std_logic_vector(7 downto 0);
    signal mulr_2_86 : std_logic_vector(7 downto 0);
    signal mulr_1_87 : std_logic_vector(7 downto 0);
    signal mulr_2_87 : std_logic_vector(7 downto 0);
    signal mulr_1_88 : std_logic_vector(7 downto 0);
    signal mulr_2_88 : std_logic_vector(7 downto 0);
    signal mulr_1_89 : std_logic_vector(7 downto 0);
    signal mulr_2_89 : std_logic_vector(7 downto 0);
    signal mulr_1_90 : std_logic_vector(7 downto 0);
    signal mulr_2_90 : std_logic_vector(7 downto 0);
    signal mulr_1_91 : std_logic_vector(7 downto 0);
    signal mulr_2_91 : std_logic_vector(7 downto 0);
    signal mulr_1_92 : std_logic_vector(7 downto 0);
    signal mulr_2_92 : std_logic_vector(7 downto 0);
    signal mulr_1_93 : std_logic_vector(7 downto 0);
    signal mulr_2_93 : std_logic_vector(7 downto 0);
    signal mulr_1_94 : std_logic_vector(7 downto 0);
    signal mulr_2_94 : std_logic_vector(7 downto 0);
    signal mulr_1_95 : std_logic_vector(7 downto 0);
    signal mulr_2_95 : std_logic_vector(7 downto 0);
    signal mulr_1_96 : std_logic_vector(7 downto 0);
    signal mulr_2_96 : std_logic_vector(7 downto 0);
    signal mulr_1_97 : std_logic_vector(7 downto 0);
    signal mulr_2_97 : std_logic_vector(7 downto 0);
    signal mulr_1_98 : std_logic_vector(7 downto 0);
    signal mulr_2_98 : std_logic_vector(7 downto 0);
    signal mulr_1_99 : std_logic_vector(7 downto 0);
    signal mulr_2_99 : std_logic_vector(7 downto 0);
    signal mulr_1_100 : std_logic_vector(7 downto 0);
    signal mulr_2_100 : std_logic_vector(7 downto 0);
    signal mulr_1_101 : std_logic_vector(7 downto 0);
    signal mulr_2_101 : std_logic_vector(7 downto 0);
    signal mulr_1_102 : std_logic_vector(7 downto 0);
    signal mulr_2_102 : std_logic_vector(7 downto 0);
    signal mulr_1_103 : std_logic_vector(7 downto 0);
    signal mulr_2_103 : std_logic_vector(7 downto 0);
    signal mulr_1_104 : std_logic_vector(7 downto 0);
    signal mulr_2_104 : std_logic_vector(7 downto 0);
    signal mulr_1_105 : std_logic_vector(7 downto 0);
    signal mulr_2_105 : std_logic_vector(7 downto 0);
    signal mulr_1_106 : std_logic_vector(7 downto 0);
    signal mulr_2_106 : std_logic_vector(7 downto 0);
    signal mulr_1_107 : std_logic_vector(7 downto 0);
    signal mulr_2_107 : std_logic_vector(7 downto 0);
    signal mulr_1_108 : std_logic_vector(7 downto 0);
    signal mulr_2_108 : std_logic_vector(7 downto 0);
    signal mulr_1_109 : std_logic_vector(7 downto 0);
    signal mulr_2_109 : std_logic_vector(7 downto 0);
    signal mulr_1_110 : std_logic_vector(7 downto 0);
    signal mulr_2_110 : std_logic_vector(7 downto 0);
    signal mulr_1_111 : std_logic_vector(7 downto 0);
    signal mulr_2_111 : std_logic_vector(7 downto 0);
    signal mulr_1_112 : std_logic_vector(7 downto 0);
    signal mulr_2_112 : std_logic_vector(7 downto 0);
    signal mulr_1_113 : std_logic_vector(7 downto 0);
    signal mulr_2_113 : std_logic_vector(7 downto 0);
    signal mulr_1_114 : std_logic_vector(7 downto 0);
    signal mulr_2_114 : std_logic_vector(7 downto 0);
    signal mulr_1_115 : std_logic_vector(7 downto 0);
    signal mulr_2_115 : std_logic_vector(7 downto 0);
    signal mulr_1_116 : std_logic_vector(7 downto 0);
    signal mulr_2_116 : std_logic_vector(7 downto 0);
    signal mulr_1_117 : std_logic_vector(7 downto 0);
    signal mulr_2_117 : std_logic_vector(7 downto 0);
    signal mulr_1_118 : std_logic_vector(7 downto 0);
    signal mulr_2_118 : std_logic_vector(7 downto 0);
    signal mulr_1_119 : std_logic_vector(7 downto 0);
    signal mulr_2_119 : std_logic_vector(7 downto 0);
    signal mulr_1_120 : std_logic_vector(7 downto 0);
    signal mulr_2_120 : std_logic_vector(7 downto 0);
    signal mulr_1_121 : std_logic_vector(7 downto 0);
    signal mulr_2_121 : std_logic_vector(7 downto 0);
    signal mulr_1_122 : std_logic_vector(7 downto 0);
    signal mulr_2_122 : std_logic_vector(7 downto 0);
    signal mulr_1_123 : std_logic_vector(7 downto 0);
    signal mulr_2_123 : std_logic_vector(7 downto 0);
    signal mulr_1_124 : std_logic_vector(7 downto 0);
    signal mulr_2_124 : std_logic_vector(7 downto 0);
    signal mulr_1_125 : std_logic_vector(7 downto 0);
    signal mulr_2_125 : std_logic_vector(7 downto 0);
    signal mulr_1_126 : std_logic_vector(7 downto 0);
    signal mulr_2_126 : std_logic_vector(7 downto 0);
    signal mulr_1_127 : std_logic_vector(7 downto 0);
    signal mulr_2_127 : std_logic_vector(7 downto 0);
    signal mulr_1_128 : std_logic_vector(7 downto 0);
    signal mulr_2_128 : std_logic_vector(7 downto 0);
    signal mulr_1_129 : std_logic_vector(7 downto 0);
    signal mulr_2_129 : std_logic_vector(7 downto 0);
    signal mulr_1_130 : std_logic_vector(7 downto 0);
    signal mulr_2_130 : std_logic_vector(7 downto 0);
    signal mulr_1_131 : std_logic_vector(7 downto 0);
    signal mulr_2_131 : std_logic_vector(7 downto 0);
    signal mulr_1_132 : std_logic_vector(7 downto 0);
    signal mulr_2_132 : std_logic_vector(7 downto 0);
    signal mulr_1_133 : std_logic_vector(7 downto 0);
    signal mulr_2_133 : std_logic_vector(7 downto 0);
    signal mulr_1_134 : std_logic_vector(7 downto 0);
    signal mulr_2_134 : std_logic_vector(7 downto 0);
    signal mulr_1_135 : std_logic_vector(7 downto 0);
    signal mulr_2_135 : std_logic_vector(7 downto 0);
    signal mulr_1_136 : std_logic_vector(7 downto 0);
    signal mulr_2_136 : std_logic_vector(7 downto 0);
    signal mulr_1_137 : std_logic_vector(7 downto 0);
    signal mulr_2_137 : std_logic_vector(7 downto 0);
    signal mulr_1_138 : std_logic_vector(7 downto 0);
    signal mulr_2_138 : std_logic_vector(7 downto 0);
    signal mulr_1_139 : std_logic_vector(7 downto 0);
    signal mulr_2_139 : std_logic_vector(7 downto 0);
    signal mulr_1_140 : std_logic_vector(7 downto 0);
    signal mulr_2_140 : std_logic_vector(7 downto 0);
    signal mulr_1_141 : std_logic_vector(7 downto 0);
    signal mulr_2_141 : std_logic_vector(7 downto 0);
    signal mulr_1_142 : std_logic_vector(7 downto 0);
    signal mulr_2_142 : std_logic_vector(7 downto 0);
    signal mulr_1_143 : std_logic_vector(7 downto 0);
    signal mulr_2_143 : std_logic_vector(7 downto 0);
    signal mulr_1_144 : std_logic_vector(7 downto 0);
    signal mulr_2_144 : std_logic_vector(7 downto 0);
    signal mulr_1_145 : std_logic_vector(7 downto 0);
    signal mulr_2_145 : std_logic_vector(7 downto 0);
    signal mulr_1_146 : std_logic_vector(7 downto 0);
    signal mulr_2_146 : std_logic_vector(7 downto 0);
    signal mulr_1_147 : std_logic_vector(7 downto 0);
    signal mulr_2_147 : std_logic_vector(7 downto 0);
    signal mulr_1_148 : std_logic_vector(7 downto 0);
    signal mulr_2_148 : std_logic_vector(7 downto 0);
    signal mulr_1_149 : std_logic_vector(7 downto 0);
    signal mulr_2_149 : std_logic_vector(7 downto 0);
    signal mulr_1_150 : std_logic_vector(7 downto 0);
    signal mulr_2_150 : std_logic_vector(7 downto 0);
    signal mulr_1_151 : std_logic_vector(7 downto 0);
    signal mulr_2_151 : std_logic_vector(7 downto 0);
    signal mulr_1_152 : std_logic_vector(7 downto 0);
    signal mulr_2_152 : std_logic_vector(7 downto 0);
    signal mulr_1_153 : std_logic_vector(7 downto 0);
    signal mulr_2_153 : std_logic_vector(7 downto 0);
    signal mulr_1_154 : std_logic_vector(7 downto 0);
    signal mulr_2_154 : std_logic_vector(7 downto 0);
    signal mulr_1_155 : std_logic_vector(7 downto 0);
    signal mulr_2_155 : std_logic_vector(7 downto 0);
    signal mulr_1_156 : std_logic_vector(7 downto 0);
    signal mulr_2_156 : std_logic_vector(7 downto 0);
    signal mulr_1_157 : std_logic_vector(7 downto 0);
    signal mulr_2_157 : std_logic_vector(7 downto 0);
    signal mulr_1_158 : std_logic_vector(7 downto 0);
    signal mulr_2_158 : std_logic_vector(7 downto 0);
    signal mulr_1_159 : std_logic_vector(7 downto 0);
    signal mulr_2_159 : std_logic_vector(7 downto 0);
    signal mulr_1_160 : std_logic_vector(7 downto 0);
    signal mulr_2_160 : std_logic_vector(7 downto 0);
    signal mulr_1_161 : std_logic_vector(7 downto 0);
    signal mulr_2_161 : std_logic_vector(7 downto 0);
    signal mulr_1_162 : std_logic_vector(7 downto 0);
    signal mulr_2_162 : std_logic_vector(7 downto 0);
    signal mulr_1_163 : std_logic_vector(7 downto 0);
    signal mulr_2_163 : std_logic_vector(7 downto 0);
    signal mulr_1_164 : std_logic_vector(7 downto 0);
    signal mulr_2_164 : std_logic_vector(7 downto 0);
    signal mulr_1_165 : std_logic_vector(7 downto 0);
    signal mulr_2_165 : std_logic_vector(7 downto 0);
    signal mulr_1_166 : std_logic_vector(7 downto 0);
    signal mulr_2_166 : std_logic_vector(7 downto 0);
    signal mulr_1_167 : std_logic_vector(7 downto 0);
    signal mulr_2_167 : std_logic_vector(7 downto 0);
    signal mulr_1_168 : std_logic_vector(7 downto 0);
    signal mulr_2_168 : std_logic_vector(7 downto 0);
    signal mulr_1_169 : std_logic_vector(7 downto 0);
    signal mulr_2_169 : std_logic_vector(7 downto 0);
    signal mulr_1_170 : std_logic_vector(7 downto 0);
    signal mulr_2_170 : std_logic_vector(7 downto 0);
    signal mulr_1_171 : std_logic_vector(7 downto 0);
    signal mulr_2_171 : std_logic_vector(7 downto 0);
    signal mulr_1_172 : std_logic_vector(7 downto 0);
    signal mulr_2_172 : std_logic_vector(7 downto 0);
    signal mulr_1_173 : std_logic_vector(7 downto 0);
    signal mulr_2_173 : std_logic_vector(7 downto 0);
    signal mulr_1_174 : std_logic_vector(7 downto 0);
    signal mulr_2_174 : std_logic_vector(7 downto 0);
    signal mulr_1_175 : std_logic_vector(7 downto 0);
    signal mulr_2_175 : std_logic_vector(7 downto 0);
    signal mulr_1_176 : std_logic_vector(7 downto 0);
    signal mulr_2_176 : std_logic_vector(7 downto 0);
    signal mulr_1_177 : std_logic_vector(7 downto 0);
    signal mulr_2_177 : std_logic_vector(7 downto 0);
    signal mulr_1_178 : std_logic_vector(7 downto 0);
    signal mulr_2_178 : std_logic_vector(7 downto 0);
    signal mulr_1_179 : std_logic_vector(7 downto 0);
    signal mulr_2_179 : std_logic_vector(7 downto 0);
    signal mulr_1_180 : std_logic_vector(7 downto 0);
    signal mulr_2_180 : std_logic_vector(7 downto 0);
    signal mulr_1_181 : std_logic_vector(7 downto 0);
    signal mulr_2_181 : std_logic_vector(7 downto 0);
    signal mulr_1_182 : std_logic_vector(7 downto 0);
    signal mulr_2_182 : std_logic_vector(7 downto 0);
    signal mulr_1_183 : std_logic_vector(7 downto 0);
    signal mulr_2_183 : std_logic_vector(7 downto 0);
    signal mulr_1_184 : std_logic_vector(7 downto 0);
    signal mulr_2_184 : std_logic_vector(7 downto 0);
    signal mulr_1_185 : std_logic_vector(7 downto 0);
    signal mulr_2_185 : std_logic_vector(7 downto 0);
    signal mulr_1_186 : std_logic_vector(7 downto 0);
    signal mulr_2_186 : std_logic_vector(7 downto 0);
    signal mulr_1_187 : std_logic_vector(7 downto 0);
    signal mulr_2_187 : std_logic_vector(7 downto 0);
    signal mulr_1_188 : std_logic_vector(7 downto 0);
    signal mulr_2_188 : std_logic_vector(7 downto 0);
    signal mulr_1_189 : std_logic_vector(7 downto 0);
    signal mulr_2_189 : std_logic_vector(7 downto 0);
    signal mulr_1_190 : std_logic_vector(7 downto 0);
    signal mulr_2_190 : std_logic_vector(7 downto 0);
    signal mulr_1_191 : std_logic_vector(7 downto 0);
    signal mulr_2_191 : std_logic_vector(7 downto 0);
    signal mulr_1_192 : std_logic_vector(7 downto 0);
    signal mulr_2_192 : std_logic_vector(7 downto 0);
    signal mulr_1_193 : std_logic_vector(7 downto 0);
    signal mulr_2_193 : std_logic_vector(7 downto 0);
    signal mulr_1_194 : std_logic_vector(7 downto 0);
    signal mulr_2_194 : std_logic_vector(7 downto 0);
    signal mulr_1_195 : std_logic_vector(7 downto 0);
    signal mulr_2_195 : std_logic_vector(7 downto 0);
    signal mulr_1_196 : std_logic_vector(7 downto 0);
    signal mulr_2_196 : std_logic_vector(7 downto 0);
    signal mulr_1_197 : std_logic_vector(7 downto 0);
    signal mulr_2_197 : std_logic_vector(7 downto 0);
    signal mulr_1_198 : std_logic_vector(7 downto 0);
    signal mulr_2_198 : std_logic_vector(7 downto 0);
    signal mulr_1_199 : std_logic_vector(7 downto 0);
    signal mulr_2_199 : std_logic_vector(7 downto 0);
    signal mulr_1_200 : std_logic_vector(7 downto 0);
    signal mulr_2_200 : std_logic_vector(7 downto 0);
    signal mulr_1_201 : std_logic_vector(7 downto 0);
    signal mulr_2_201 : std_logic_vector(7 downto 0);
    signal mulr_1_202 : std_logic_vector(7 downto 0);
    signal mulr_2_202 : std_logic_vector(7 downto 0);
    signal mulr_1_203 : std_logic_vector(7 downto 0);
    signal mulr_2_203 : std_logic_vector(7 downto 0);
    signal mulr_1_204 : std_logic_vector(7 downto 0);
    signal mulr_2_204 : std_logic_vector(7 downto 0);
    signal mulr_1_205 : std_logic_vector(7 downto 0);
    signal mulr_2_205 : std_logic_vector(7 downto 0);
    signal mulr_1_206 : std_logic_vector(7 downto 0);
    signal mulr_2_206 : std_logic_vector(7 downto 0);
    signal mulr_1_207 : std_logic_vector(7 downto 0);
    signal mulr_2_207 : std_logic_vector(7 downto 0);
    signal mulr_1_208 : std_logic_vector(7 downto 0);
    signal mulr_2_208 : std_logic_vector(7 downto 0);
    signal mulr_1_209 : std_logic_vector(7 downto 0);
    signal mulr_2_209 : std_logic_vector(7 downto 0);
    signal mulr_1_210 : std_logic_vector(7 downto 0);
    signal mulr_2_210 : std_logic_vector(7 downto 0);
    signal mulr_1_211 : std_logic_vector(7 downto 0);
    signal mulr_2_211 : std_logic_vector(7 downto 0);
    signal mulr_1_212 : std_logic_vector(7 downto 0);
    signal mulr_2_212 : std_logic_vector(7 downto 0);
    signal mulr_1_213 : std_logic_vector(7 downto 0);
    signal mulr_2_213 : std_logic_vector(7 downto 0);
    signal mulr_1_214 : std_logic_vector(7 downto 0);
    signal mulr_2_214 : std_logic_vector(7 downto 0);
    signal mulr_1_215 : std_logic_vector(7 downto 0);
    signal mulr_2_215 : std_logic_vector(7 downto 0);
    signal mulr_1_216 : std_logic_vector(7 downto 0);
    signal mulr_2_216 : std_logic_vector(7 downto 0);
    signal mulr_1_217 : std_logic_vector(7 downto 0);
    signal mulr_2_217 : std_logic_vector(7 downto 0);
    signal mulr_1_218 : std_logic_vector(7 downto 0);
    signal mulr_2_218 : std_logic_vector(7 downto 0);
    signal mulr_1_219 : std_logic_vector(7 downto 0);
    signal mulr_2_219 : std_logic_vector(7 downto 0);
    signal mulr_1_220 : std_logic_vector(7 downto 0);
    signal mulr_2_220 : std_logic_vector(7 downto 0);
    signal mulr_1_221 : std_logic_vector(7 downto 0);
    signal mulr_2_221 : std_logic_vector(7 downto 0);
    signal mulr_1_222 : std_logic_vector(7 downto 0);
    signal mulr_2_222 : std_logic_vector(7 downto 0);
    signal mulr_1_223 : std_logic_vector(7 downto 0);
    signal mulr_2_223 : std_logic_vector(7 downto 0);
    signal mulr_1_224 : std_logic_vector(7 downto 0);
    signal mulr_2_224 : std_logic_vector(7 downto 0);
    signal mulr_1_225 : std_logic_vector(7 downto 0);
    signal mulr_2_225 : std_logic_vector(7 downto 0);
    signal mulr_1_226 : std_logic_vector(7 downto 0);
    signal mulr_2_226 : std_logic_vector(7 downto 0);
    signal mulr_1_227 : std_logic_vector(7 downto 0);
    signal mulr_2_227 : std_logic_vector(7 downto 0);
    signal mulr_1_228 : std_logic_vector(7 downto 0);
    signal mulr_2_228 : std_logic_vector(7 downto 0);
    signal mulr_1_229 : std_logic_vector(7 downto 0);
    signal mulr_2_229 : std_logic_vector(7 downto 0);
    signal mulr_1_230 : std_logic_vector(7 downto 0);
    signal mulr_2_230 : std_logic_vector(7 downto 0);
    signal mulr_1_231 : std_logic_vector(7 downto 0);
    signal mulr_2_231 : std_logic_vector(7 downto 0);
    signal mulr_1_232 : std_logic_vector(7 downto 0);
    signal mulr_2_232 : std_logic_vector(7 downto 0);
    signal mulr_1_233 : std_logic_vector(7 downto 0);
    signal mulr_2_233 : std_logic_vector(7 downto 0);
    signal mulr_1_234 : std_logic_vector(7 downto 0);
    signal mulr_2_234 : std_logic_vector(7 downto 0);
    signal mulr_1_235 : std_logic_vector(7 downto 0);
    signal mulr_2_235 : std_logic_vector(7 downto 0);
    signal mulr_1_236 : std_logic_vector(7 downto 0);
    signal mulr_2_236 : std_logic_vector(7 downto 0);
    signal mulr_1_237 : std_logic_vector(7 downto 0);
    signal mulr_2_237 : std_logic_vector(7 downto 0);
    signal mulr_1_238 : std_logic_vector(7 downto 0);
    signal mulr_2_238 : std_logic_vector(7 downto 0);
    signal mulr_1_239 : std_logic_vector(7 downto 0);
    signal mulr_2_239 : std_logic_vector(7 downto 0);
    signal mulr_1_240 : std_logic_vector(7 downto 0);
    signal mulr_2_240 : std_logic_vector(7 downto 0);
    signal mulr_1_241 : std_logic_vector(7 downto 0);
    signal mulr_2_241 : std_logic_vector(7 downto 0);
    signal mulr_1_242 : std_logic_vector(7 downto 0);
    signal mulr_2_242 : std_logic_vector(7 downto 0);
    signal mulr_1_243 : std_logic_vector(7 downto 0);
    signal mulr_2_243 : std_logic_vector(7 downto 0);
    signal mulr_1_244 : std_logic_vector(7 downto 0);
    signal mulr_2_244 : std_logic_vector(7 downto 0);
    signal mulr_1_245 : std_logic_vector(7 downto 0);
    signal mulr_2_245 : std_logic_vector(7 downto 0);
    signal mulr_1_246 : std_logic_vector(7 downto 0);
    signal mulr_2_246 : std_logic_vector(7 downto 0);
    signal mulr_1_247 : std_logic_vector(7 downto 0);
    signal mulr_2_247 : std_logic_vector(7 downto 0);
    signal mulr_1_248 : std_logic_vector(7 downto 0);
    signal mulr_2_248 : std_logic_vector(7 downto 0);
    signal mulr_1_249 : std_logic_vector(7 downto 0);
    signal mulr_2_249 : std_logic_vector(7 downto 0);
    signal mulr_1_250 : std_logic_vector(7 downto 0);
    signal mulr_2_250 : std_logic_vector(7 downto 0);
    signal mulr_1_251 : std_logic_vector(7 downto 0);
    signal mulr_2_251 : std_logic_vector(7 downto 0);
    signal mulr_1_252 : std_logic_vector(7 downto 0);
    signal mulr_2_252 : std_logic_vector(7 downto 0);
    signal mulr_1_253 : std_logic_vector(7 downto 0);
    signal mulr_2_253 : std_logic_vector(7 downto 0);
    signal mulr_1_254 : std_logic_vector(7 downto 0);
    signal mulr_2_254 : std_logic_vector(7 downto 0);
    signal mulr_1_255 : std_logic_vector(7 downto 0);
    signal mulr_2_255 : std_logic_vector(7 downto 0);
    signal sumr_1 : std_logic_vector(7 downto 0);
    signal sumr_2 : std_logic_vector(7 downto 0);
    signal sumr_3 : std_logic_vector(7 downto 0);
    signal sumr_4 : std_logic_vector(7 downto 0);
    signal sumr_5 : std_logic_vector(7 downto 0);
    signal sumr_6 : std_logic_vector(7 downto 0);
    signal sumr_7 : std_logic_vector(7 downto 0);
    signal sumr_8 : std_logic_vector(7 downto 0);
    signal sumr_9 : std_logic_vector(7 downto 0);
    signal sumr_10 : std_logic_vector(7 downto 0);
    signal sumr_11 : std_logic_vector(7 downto 0);
    signal sumr_12 : std_logic_vector(7 downto 0);
    signal sumr_13 : std_logic_vector(7 downto 0);
    signal sumr_14 : std_logic_vector(7 downto 0);
    signal sumr_15 : std_logic_vector(7 downto 0);
    signal sumr_16 : std_logic_vector(7 downto 0);
    signal sumr_17 : std_logic_vector(7 downto 0);
    signal sumr_18 : std_logic_vector(7 downto 0);
    signal sumr_19 : std_logic_vector(7 downto 0);
    signal sumr_20 : std_logic_vector(7 downto 0);
    signal sumr_21 : std_logic_vector(7 downto 0);
    signal sumr_22 : std_logic_vector(7 downto 0);
    signal sumr_23 : std_logic_vector(7 downto 0);
    signal sumr_24 : std_logic_vector(7 downto 0);
    signal sumr_25 : std_logic_vector(7 downto 0);
    signal sumr_26 : std_logic_vector(7 downto 0);
    signal sumr_27 : std_logic_vector(7 downto 0);
    signal sumr_28 : std_logic_vector(7 downto 0);
    signal sumr_29 : std_logic_vector(7 downto 0);
    signal sumr_30 : std_logic_vector(7 downto 0);
    signal sumr_31 : std_logic_vector(7 downto 0);
    signal sumr_32 : std_logic_vector(7 downto 0);
    signal sumr_33 : std_logic_vector(7 downto 0);
    signal sumr_34 : std_logic_vector(7 downto 0);
    signal sumr_35 : std_logic_vector(7 downto 0);
    signal sumr_36 : std_logic_vector(7 downto 0);
    signal sumr_37 : std_logic_vector(7 downto 0);
    signal sumr_38 : std_logic_vector(7 downto 0);
    signal sumr_39 : std_logic_vector(7 downto 0);
    signal sumr_40 : std_logic_vector(7 downto 0);
    signal sumr_41 : std_logic_vector(7 downto 0);
    signal sumr_42 : std_logic_vector(7 downto 0);
    signal sumr_43 : std_logic_vector(7 downto 0);
    signal sumr_44 : std_logic_vector(7 downto 0);
    signal sumr_45 : std_logic_vector(7 downto 0);
    signal sumr_46 : std_logic_vector(7 downto 0);
    signal sumr_47 : std_logic_vector(7 downto 0);
    signal sumr_48 : std_logic_vector(7 downto 0);
    signal sumr_49 : std_logic_vector(7 downto 0);
    signal sumr_50 : std_logic_vector(7 downto 0);
    signal sumr_51 : std_logic_vector(7 downto 0);
    signal sumr_52 : std_logic_vector(7 downto 0);
    signal sumr_53 : std_logic_vector(7 downto 0);
    signal sumr_54 : std_logic_vector(7 downto 0);
    signal sumr_55 : std_logic_vector(7 downto 0);
    signal sumr_56 : std_logic_vector(7 downto 0);
    signal sumr_57 : std_logic_vector(7 downto 0);
    signal sumr_58 : std_logic_vector(7 downto 0);
    signal sumr_59 : std_logic_vector(7 downto 0);
    signal sumr_60 : std_logic_vector(7 downto 0);
    signal sumr_61 : std_logic_vector(7 downto 0);
    signal sumr_62 : std_logic_vector(7 downto 0);
    signal sumr_63 : std_logic_vector(7 downto 0);
    signal sumr_64 : std_logic_vector(7 downto 0);
    signal sumr_65 : std_logic_vector(7 downto 0);
    signal sumr_66 : std_logic_vector(7 downto 0);
    signal sumr_67 : std_logic_vector(7 downto 0);
    signal sumr_68 : std_logic_vector(7 downto 0);
    signal sumr_69 : std_logic_vector(7 downto 0);
    signal sumr_70 : std_logic_vector(7 downto 0);
    signal sumr_71 : std_logic_vector(7 downto 0);
    signal sumr_72 : std_logic_vector(7 downto 0);
    signal sumr_73 : std_logic_vector(7 downto 0);
    signal sumr_74 : std_logic_vector(7 downto 0);
    signal sumr_75 : std_logic_vector(7 downto 0);
    signal sumr_76 : std_logic_vector(7 downto 0);
    signal sumr_77 : std_logic_vector(7 downto 0);
    signal sumr_78 : std_logic_vector(7 downto 0);
    signal sumr_79 : std_logic_vector(7 downto 0);
    signal sumr_80 : std_logic_vector(7 downto 0);
    signal sumr_81 : std_logic_vector(7 downto 0);
    signal sumr_82 : std_logic_vector(7 downto 0);
    signal sumr_83 : std_logic_vector(7 downto 0);
    signal sumr_84 : std_logic_vector(7 downto 0);
    signal sumr_85 : std_logic_vector(7 downto 0);
    signal sumr_86 : std_logic_vector(7 downto 0);
    signal sumr_87 : std_logic_vector(7 downto 0);
    signal sumr_88 : std_logic_vector(7 downto 0);
    signal sumr_89 : std_logic_vector(7 downto 0);
    signal sumr_90 : std_logic_vector(7 downto 0);
    signal sumr_91 : std_logic_vector(7 downto 0);
    signal sumr_92 : std_logic_vector(7 downto 0);
    signal sumr_93 : std_logic_vector(7 downto 0);
    signal sumr_94 : std_logic_vector(7 downto 0);
    signal sumr_95 : std_logic_vector(7 downto 0);
    signal sumr_96 : std_logic_vector(7 downto 0);
    signal sumr_97 : std_logic_vector(7 downto 0);
    signal sumr_98 : std_logic_vector(7 downto 0);
    signal sumr_99 : std_logic_vector(7 downto 0);
    signal sumr_100 : std_logic_vector(7 downto 0);
    signal sumr_101 : std_logic_vector(7 downto 0);
    signal sumr_102 : std_logic_vector(7 downto 0);
    signal sumr_103 : std_logic_vector(7 downto 0);
    signal sumr_104 : std_logic_vector(7 downto 0);
    signal sumr_105 : std_logic_vector(7 downto 0);
    signal sumr_106 : std_logic_vector(7 downto 0);
    signal sumr_107 : std_logic_vector(7 downto 0);
    signal sumr_108 : std_logic_vector(7 downto 0);
    signal sumr_109 : std_logic_vector(7 downto 0);
    signal sumr_110 : std_logic_vector(7 downto 0);
    signal sumr_111 : std_logic_vector(7 downto 0);
    signal sumr_112 : std_logic_vector(7 downto 0);
    signal sumr_113 : std_logic_vector(7 downto 0);
    signal sumr_114 : std_logic_vector(7 downto 0);
    signal sumr_115 : std_logic_vector(7 downto 0);
    signal sumr_116 : std_logic_vector(7 downto 0);
    signal sumr_117 : std_logic_vector(7 downto 0);
    signal sumr_118 : std_logic_vector(7 downto 0);
    signal sumr_119 : std_logic_vector(7 downto 0);
    signal sumr_120 : std_logic_vector(7 downto 0);
    signal sumr_121 : std_logic_vector(7 downto 0);
    signal sumr_122 : std_logic_vector(7 downto 0);
    signal sumr_123 : std_logic_vector(7 downto 0);
    signal sumr_124 : std_logic_vector(7 downto 0);
    signal sumr_125 : std_logic_vector(7 downto 0);
    signal sumr_126 : std_logic_vector(7 downto 0);
    signal sumr_127 : std_logic_vector(7 downto 0);
    signal sumr_128 : std_logic_vector(7 downto 0);
    signal sumr_129 : std_logic_vector(7 downto 0);
    signal sumr_130 : std_logic_vector(7 downto 0);
    signal sumr_131 : std_logic_vector(7 downto 0);
    signal sumr_132 : std_logic_vector(7 downto 0);
    signal sumr_133 : std_logic_vector(7 downto 0);
    signal sumr_134 : std_logic_vector(7 downto 0);
    signal sumr_135 : std_logic_vector(7 downto 0);
    signal sumr_136 : std_logic_vector(7 downto 0);
    signal sumr_137 : std_logic_vector(7 downto 0);
    signal sumr_138 : std_logic_vector(7 downto 0);
    signal sumr_139 : std_logic_vector(7 downto 0);
    signal sumr_140 : std_logic_vector(7 downto 0);
    signal sumr_141 : std_logic_vector(7 downto 0);
    signal sumr_142 : std_logic_vector(7 downto 0);
    signal sumr_143 : std_logic_vector(7 downto 0);
    signal sumr_144 : std_logic_vector(7 downto 0);
    signal sumr_145 : std_logic_vector(7 downto 0);
    signal sumr_146 : std_logic_vector(7 downto 0);
    signal sumr_147 : std_logic_vector(7 downto 0);
    signal sumr_148 : std_logic_vector(7 downto 0);
    signal sumr_149 : std_logic_vector(7 downto 0);
    signal sumr_150 : std_logic_vector(7 downto 0);
    signal sumr_151 : std_logic_vector(7 downto 0);
    signal sumr_152 : std_logic_vector(7 downto 0);
    signal sumr_153 : std_logic_vector(7 downto 0);
    signal sumr_154 : std_logic_vector(7 downto 0);
    signal sumr_155 : std_logic_vector(7 downto 0);
    signal sumr_156 : std_logic_vector(7 downto 0);
    signal sumr_157 : std_logic_vector(7 downto 0);
    signal sumr_158 : std_logic_vector(7 downto 0);
    signal sumr_159 : std_logic_vector(7 downto 0);
    signal sumr_160 : std_logic_vector(7 downto 0);
    signal sumr_161 : std_logic_vector(7 downto 0);
    signal sumr_162 : std_logic_vector(7 downto 0);
    signal sumr_163 : std_logic_vector(7 downto 0);
    signal sumr_164 : std_logic_vector(7 downto 0);
    signal sumr_165 : std_logic_vector(7 downto 0);
    signal sumr_166 : std_logic_vector(7 downto 0);
    signal sumr_167 : std_logic_vector(7 downto 0);
    signal sumr_168 : std_logic_vector(7 downto 0);
    signal sumr_169 : std_logic_vector(7 downto 0);
    signal sumr_170 : std_logic_vector(7 downto 0);
    signal sumr_171 : std_logic_vector(7 downto 0);
    signal sumr_172 : std_logic_vector(7 downto 0);
    signal sumr_173 : std_logic_vector(7 downto 0);
    signal sumr_174 : std_logic_vector(7 downto 0);
    signal sumr_175 : std_logic_vector(7 downto 0);
    signal sumr_176 : std_logic_vector(7 downto 0);
    signal sumr_177 : std_logic_vector(7 downto 0);
    signal sumr_178 : std_logic_vector(7 downto 0);
    signal sumr_179 : std_logic_vector(7 downto 0);
    signal sumr_180 : std_logic_vector(7 downto 0);
    signal sumr_181 : std_logic_vector(7 downto 0);
    signal sumr_182 : std_logic_vector(7 downto 0);
    signal sumr_183 : std_logic_vector(7 downto 0);
    signal sumr_184 : std_logic_vector(7 downto 0);
    signal sumr_185 : std_logic_vector(7 downto 0);
    signal sumr_186 : std_logic_vector(7 downto 0);
    signal sumr_187 : std_logic_vector(7 downto 0);
    signal sumr_188 : std_logic_vector(7 downto 0);
    signal sumr_189 : std_logic_vector(7 downto 0);
    signal sumr_190 : std_logic_vector(7 downto 0);
    signal sumr_191 : std_logic_vector(7 downto 0);
    signal sumr_192 : std_logic_vector(7 downto 0);
    signal sumr_193 : std_logic_vector(7 downto 0);
    signal sumr_194 : std_logic_vector(7 downto 0);
    signal sumr_195 : std_logic_vector(7 downto 0);
    signal sumr_196 : std_logic_vector(7 downto 0);
    signal sumr_197 : std_logic_vector(7 downto 0);
    signal sumr_198 : std_logic_vector(7 downto 0);
    signal sumr_199 : std_logic_vector(7 downto 0);
    signal sumr_200 : std_logic_vector(7 downto 0);
    signal sumr_201 : std_logic_vector(7 downto 0);
    signal sumr_202 : std_logic_vector(7 downto 0);
    signal sumr_203 : std_logic_vector(7 downto 0);
    signal sumr_204 : std_logic_vector(7 downto 0);
    signal sumr_205 : std_logic_vector(7 downto 0);
    signal sumr_206 : std_logic_vector(7 downto 0);
    signal sumr_207 : std_logic_vector(7 downto 0);
    signal sumr_208 : std_logic_vector(7 downto 0);
    signal sumr_209 : std_logic_vector(7 downto 0);
    signal sumr_210 : std_logic_vector(7 downto 0);
    signal sumr_211 : std_logic_vector(7 downto 0);
    signal sumr_212 : std_logic_vector(7 downto 0);
    signal sumr_213 : std_logic_vector(7 downto 0);
    signal sumr_214 : std_logic_vector(7 downto 0);
    signal sumr_215 : std_logic_vector(7 downto 0);
    signal sumr_216 : std_logic_vector(7 downto 0);
    signal sumr_217 : std_logic_vector(7 downto 0);
    signal sumr_218 : std_logic_vector(7 downto 0);
    signal sumr_219 : std_logic_vector(7 downto 0);
    signal sumr_220 : std_logic_vector(7 downto 0);
    signal sumr_221 : std_logic_vector(7 downto 0);
    signal sumr_222 : std_logic_vector(7 downto 0);
    signal sumr_223 : std_logic_vector(7 downto 0);
    signal sumr_224 : std_logic_vector(7 downto 0);
    signal sumr_225 : std_logic_vector(7 downto 0);
    signal sumr_226 : std_logic_vector(7 downto 0);
    signal sumr_227 : std_logic_vector(7 downto 0);
    signal sumr_228 : std_logic_vector(7 downto 0);
    signal sumr_229 : std_logic_vector(7 downto 0);
    signal sumr_230 : std_logic_vector(7 downto 0);
    signal sumr_231 : std_logic_vector(7 downto 0);
    signal sumr_232 : std_logic_vector(7 downto 0);
    signal sumr_233 : std_logic_vector(7 downto 0);
    signal sumr_234 : std_logic_vector(7 downto 0);
    signal sumr_235 : std_logic_vector(7 downto 0);
    signal sumr_236 : std_logic_vector(7 downto 0);
    signal sumr_237 : std_logic_vector(7 downto 0);
    signal sumr_238 : std_logic_vector(7 downto 0);
    signal sumr_239 : std_logic_vector(7 downto 0);
    signal sumr_240 : std_logic_vector(7 downto 0);
    signal sumr_241 : std_logic_vector(7 downto 0);
    signal sumr_242 : std_logic_vector(7 downto 0);
    signal sumr_243 : std_logic_vector(7 downto 0);
    signal sumr_244 : std_logic_vector(7 downto 0);
    signal sumr_245 : std_logic_vector(7 downto 0);
    signal sumr_246 : std_logic_vector(7 downto 0);
    signal sumr_247 : std_logic_vector(7 downto 0);
    signal sumr_248 : std_logic_vector(7 downto 0);
    signal sumr_249 : std_logic_vector(7 downto 0);
    signal sumr_250 : std_logic_vector(7 downto 0);
    signal sumr_251 : std_logic_vector(7 downto 0);
    signal sumr_252 : std_logic_vector(7 downto 0);
    signal sumr_253 : std_logic_vector(7 downto 0);
    signal sumr_254 : std_logic_vector(7 downto 0);
    signal sumr_255 : std_logic_vector(7 downto 0);
begin

mulr_1_1<=a_1;
mulc_2_1 : entity work.gfmul
port map(
a=>a_2,
b=>"00000010",
X=>mulr_2_1);

mulr_1_2<=a_1;
mulc_2_2 : entity work.gfmul
port map(
a=>a_2,
b=>"00000100",
X=>mulr_2_2);

mulr_1_3<=a_1;
mulc_2_3 : entity work.gfmul
port map(
a=>a_2,
b=>"00001000",
X=>mulr_2_3);

mulr_1_4<=a_1;
mulc_2_4 : entity work.gfmul
port map(
a=>a_2,
b=>"00010000",
X=>mulr_2_4);

mulr_1_5<=a_1;
mulc_2_5 : entity work.gfmul
port map(
a=>a_2,
b=>"00100000",
X=>mulr_2_5);

mulr_1_6<=a_1;
mulc_2_6 : entity work.gfmul
port map(
a=>a_2,
b=>"01000000",
X=>mulr_2_6);

mulr_1_7<=a_1;
mulc_2_7 : entity work.gfmul
port map(
a=>a_2,
b=>"10000000",
X=>mulr_2_7);

mulr_1_8<=a_1;
mulc_2_8 : entity work.gfmul
port map(
a=>a_2,
b=>"00011101",
X=>mulr_2_8);

mulr_1_9<=a_1;
mulc_2_9 : entity work.gfmul
port map(
a=>a_2,
b=>"00111010",
X=>mulr_2_9);

mulr_1_10<=a_1;
mulc_2_10 : entity work.gfmul
port map(
a=>a_2,
b=>"01110100",
X=>mulr_2_10);

mulr_1_11<=a_1;
mulc_2_11 : entity work.gfmul
port map(
a=>a_2,
b=>"11101000",
X=>mulr_2_11);

mulr_1_12<=a_1;
mulc_2_12 : entity work.gfmul
port map(
a=>a_2,
b=>"11001101",
X=>mulr_2_12);

mulr_1_13<=a_1;
mulc_2_13 : entity work.gfmul
port map(
a=>a_2,
b=>"10000111",
X=>mulr_2_13);

mulr_1_14<=a_1;
mulc_2_14 : entity work.gfmul
port map(
a=>a_2,
b=>"00010011",
X=>mulr_2_14);

mulr_1_15<=a_1;
mulc_2_15 : entity work.gfmul
port map(
a=>a_2,
b=>"00100110",
X=>mulr_2_15);

mulr_1_16<=a_1;
mulc_2_16 : entity work.gfmul
port map(
a=>a_2,
b=>"01001100",
X=>mulr_2_16);

mulr_1_17<=a_1;
mulc_2_17 : entity work.gfmul
port map(
a=>a_2,
b=>"10011000",
X=>mulr_2_17);

mulr_1_18<=a_1;
mulc_2_18 : entity work.gfmul
port map(
a=>a_2,
b=>"00101101",
X=>mulr_2_18);

mulr_1_19<=a_1;
mulc_2_19 : entity work.gfmul
port map(
a=>a_2,
b=>"01011010",
X=>mulr_2_19);

mulr_1_20<=a_1;
mulc_2_20 : entity work.gfmul
port map(
a=>a_2,
b=>"10110100",
X=>mulr_2_20);

mulr_1_21<=a_1;
mulc_2_21 : entity work.gfmul
port map(
a=>a_2,
b=>"01110101",
X=>mulr_2_21);

mulr_1_22<=a_1;
mulc_2_22 : entity work.gfmul
port map(
a=>a_2,
b=>"11101010",
X=>mulr_2_22);

mulr_1_23<=a_1;
mulc_2_23 : entity work.gfmul
port map(
a=>a_2,
b=>"11001001",
X=>mulr_2_23);

mulr_1_24<=a_1;
mulc_2_24 : entity work.gfmul
port map(
a=>a_2,
b=>"10001111",
X=>mulr_2_24);

mulr_1_25<=a_1;
mulc_2_25 : entity work.gfmul
port map(
a=>a_2,
b=>"00000011",
X=>mulr_2_25);

mulr_1_26<=a_1;
mulc_2_26 : entity work.gfmul
port map(
a=>a_2,
b=>"00000110",
X=>mulr_2_26);

mulr_1_27<=a_1;
mulc_2_27 : entity work.gfmul
port map(
a=>a_2,
b=>"00001100",
X=>mulr_2_27);

mulr_1_28<=a_1;
mulc_2_28 : entity work.gfmul
port map(
a=>a_2,
b=>"00011000",
X=>mulr_2_28);

mulr_1_29<=a_1;
mulc_2_29 : entity work.gfmul
port map(
a=>a_2,
b=>"00110000",
X=>mulr_2_29);

mulr_1_30<=a_1;
mulc_2_30 : entity work.gfmul
port map(
a=>a_2,
b=>"01100000",
X=>mulr_2_30);

mulr_1_31<=a_1;
mulc_2_31 : entity work.gfmul
port map(
a=>a_2,
b=>"11000000",
X=>mulr_2_31);

mulr_1_32<=a_1;
mulc_2_32 : entity work.gfmul
port map(
a=>a_2,
b=>"10011101",
X=>mulr_2_32);

mulr_1_33<=a_1;
mulc_2_33 : entity work.gfmul
port map(
a=>a_2,
b=>"00100111",
X=>mulr_2_33);

mulr_1_34<=a_1;
mulc_2_34 : entity work.gfmul
port map(
a=>a_2,
b=>"01001110",
X=>mulr_2_34);

mulr_1_35<=a_1;
mulc_2_35 : entity work.gfmul
port map(
a=>a_2,
b=>"10011100",
X=>mulr_2_35);

mulr_1_36<=a_1;
mulc_2_36 : entity work.gfmul
port map(
a=>a_2,
b=>"00100101",
X=>mulr_2_36);

mulr_1_37<=a_1;
mulc_2_37 : entity work.gfmul
port map(
a=>a_2,
b=>"01001010",
X=>mulr_2_37);

mulr_1_38<=a_1;
mulc_2_38 : entity work.gfmul
port map(
a=>a_2,
b=>"10010100",
X=>mulr_2_38);

mulr_1_39<=a_1;
mulc_2_39 : entity work.gfmul
port map(
a=>a_2,
b=>"00110101",
X=>mulr_2_39);

mulr_1_40<=a_1;
mulc_2_40 : entity work.gfmul
port map(
a=>a_2,
b=>"01101010",
X=>mulr_2_40);

mulr_1_41<=a_1;
mulc_2_41 : entity work.gfmul
port map(
a=>a_2,
b=>"11010100",
X=>mulr_2_41);

mulr_1_42<=a_1;
mulc_2_42 : entity work.gfmul
port map(
a=>a_2,
b=>"10110101",
X=>mulr_2_42);

mulr_1_43<=a_1;
mulc_2_43 : entity work.gfmul
port map(
a=>a_2,
b=>"01110111",
X=>mulr_2_43);

mulr_1_44<=a_1;
mulc_2_44 : entity work.gfmul
port map(
a=>a_2,
b=>"11101110",
X=>mulr_2_44);

mulr_1_45<=a_1;
mulc_2_45 : entity work.gfmul
port map(
a=>a_2,
b=>"11000001",
X=>mulr_2_45);

mulr_1_46<=a_1;
mulc_2_46 : entity work.gfmul
port map(
a=>a_2,
b=>"10011111",
X=>mulr_2_46);

mulr_1_47<=a_1;
mulc_2_47 : entity work.gfmul
port map(
a=>a_2,
b=>"00100011",
X=>mulr_2_47);

mulr_1_48<=a_1;
mulc_2_48 : entity work.gfmul
port map(
a=>a_2,
b=>"01000110",
X=>mulr_2_48);

mulr_1_49<=a_1;
mulc_2_49 : entity work.gfmul
port map(
a=>a_2,
b=>"10001100",
X=>mulr_2_49);

mulr_1_50<=a_1;
mulc_2_50 : entity work.gfmul
port map(
a=>a_2,
b=>"00000101",
X=>mulr_2_50);

mulr_1_51<=a_1;
mulc_2_51 : entity work.gfmul
port map(
a=>a_2,
b=>"00001010",
X=>mulr_2_51);

mulr_1_52<=a_1;
mulc_2_52 : entity work.gfmul
port map(
a=>a_2,
b=>"00010100",
X=>mulr_2_52);

mulr_1_53<=a_1;
mulc_2_53 : entity work.gfmul
port map(
a=>a_2,
b=>"00101000",
X=>mulr_2_53);

mulr_1_54<=a_1;
mulc_2_54 : entity work.gfmul
port map(
a=>a_2,
b=>"01010000",
X=>mulr_2_54);

mulr_1_55<=a_1;
mulc_2_55 : entity work.gfmul
port map(
a=>a_2,
b=>"10100000",
X=>mulr_2_55);

mulr_1_56<=a_1;
mulc_2_56 : entity work.gfmul
port map(
a=>a_2,
b=>"01011101",
X=>mulr_2_56);

mulr_1_57<=a_1;
mulc_2_57 : entity work.gfmul
port map(
a=>a_2,
b=>"10111010",
X=>mulr_2_57);

mulr_1_58<=a_1;
mulc_2_58 : entity work.gfmul
port map(
a=>a_2,
b=>"01101001",
X=>mulr_2_58);

mulr_1_59<=a_1;
mulc_2_59 : entity work.gfmul
port map(
a=>a_2,
b=>"11010010",
X=>mulr_2_59);

mulr_1_60<=a_1;
mulc_2_60 : entity work.gfmul
port map(
a=>a_2,
b=>"10111001",
X=>mulr_2_60);

mulr_1_61<=a_1;
mulc_2_61 : entity work.gfmul
port map(
a=>a_2,
b=>"01101111",
X=>mulr_2_61);

mulr_1_62<=a_1;
mulc_2_62 : entity work.gfmul
port map(
a=>a_2,
b=>"11011110",
X=>mulr_2_62);

mulr_1_63<=a_1;
mulc_2_63 : entity work.gfmul
port map(
a=>a_2,
b=>"10100001",
X=>mulr_2_63);

mulr_1_64<=a_1;
mulc_2_64 : entity work.gfmul
port map(
a=>a_2,
b=>"01011111",
X=>mulr_2_64);

mulr_1_65<=a_1;
mulc_2_65 : entity work.gfmul
port map(
a=>a_2,
b=>"10111110",
X=>mulr_2_65);

mulr_1_66<=a_1;
mulc_2_66 : entity work.gfmul
port map(
a=>a_2,
b=>"01100001",
X=>mulr_2_66);

mulr_1_67<=a_1;
mulc_2_67 : entity work.gfmul
port map(
a=>a_2,
b=>"11000010",
X=>mulr_2_67);

mulr_1_68<=a_1;
mulc_2_68 : entity work.gfmul
port map(
a=>a_2,
b=>"10011001",
X=>mulr_2_68);

mulr_1_69<=a_1;
mulc_2_69 : entity work.gfmul
port map(
a=>a_2,
b=>"00101111",
X=>mulr_2_69);

mulr_1_70<=a_1;
mulc_2_70 : entity work.gfmul
port map(
a=>a_2,
b=>"01011110",
X=>mulr_2_70);

mulr_1_71<=a_1;
mulc_2_71 : entity work.gfmul
port map(
a=>a_2,
b=>"10111100",
X=>mulr_2_71);

mulr_1_72<=a_1;
mulc_2_72 : entity work.gfmul
port map(
a=>a_2,
b=>"01100101",
X=>mulr_2_72);

mulr_1_73<=a_1;
mulc_2_73 : entity work.gfmul
port map(
a=>a_2,
b=>"11001010",
X=>mulr_2_73);

mulr_1_74<=a_1;
mulc_2_74 : entity work.gfmul
port map(
a=>a_2,
b=>"10001001",
X=>mulr_2_74);

mulr_1_75<=a_1;
mulc_2_75 : entity work.gfmul
port map(
a=>a_2,
b=>"00001111",
X=>mulr_2_75);

mulr_1_76<=a_1;
mulc_2_76 : entity work.gfmul
port map(
a=>a_2,
b=>"00011110",
X=>mulr_2_76);

mulr_1_77<=a_1;
mulc_2_77 : entity work.gfmul
port map(
a=>a_2,
b=>"00111100",
X=>mulr_2_77);

mulr_1_78<=a_1;
mulc_2_78 : entity work.gfmul
port map(
a=>a_2,
b=>"01111000",
X=>mulr_2_78);

mulr_1_79<=a_1;
mulc_2_79 : entity work.gfmul
port map(
a=>a_2,
b=>"11110000",
X=>mulr_2_79);

mulr_1_80<=a_1;
mulc_2_80 : entity work.gfmul
port map(
a=>a_2,
b=>"11111101",
X=>mulr_2_80);

mulr_1_81<=a_1;
mulc_2_81 : entity work.gfmul
port map(
a=>a_2,
b=>"11100111",
X=>mulr_2_81);

mulr_1_82<=a_1;
mulc_2_82 : entity work.gfmul
port map(
a=>a_2,
b=>"11010011",
X=>mulr_2_82);

mulr_1_83<=a_1;
mulc_2_83 : entity work.gfmul
port map(
a=>a_2,
b=>"10111011",
X=>mulr_2_83);

mulr_1_84<=a_1;
mulc_2_84 : entity work.gfmul
port map(
a=>a_2,
b=>"01101011",
X=>mulr_2_84);

mulr_1_85<=a_1;
mulc_2_85 : entity work.gfmul
port map(
a=>a_2,
b=>"11010110",
X=>mulr_2_85);

mulr_1_86<=a_1;
mulc_2_86 : entity work.gfmul
port map(
a=>a_2,
b=>"10110001",
X=>mulr_2_86);

mulr_1_87<=a_1;
mulc_2_87 : entity work.gfmul
port map(
a=>a_2,
b=>"01111111",
X=>mulr_2_87);

mulr_1_88<=a_1;
mulc_2_88 : entity work.gfmul
port map(
a=>a_2,
b=>"11111110",
X=>mulr_2_88);

mulr_1_89<=a_1;
mulc_2_89 : entity work.gfmul
port map(
a=>a_2,
b=>"11100001",
X=>mulr_2_89);

mulr_1_90<=a_1;
mulc_2_90 : entity work.gfmul
port map(
a=>a_2,
b=>"11011111",
X=>mulr_2_90);

mulr_1_91<=a_1;
mulc_2_91 : entity work.gfmul
port map(
a=>a_2,
b=>"10100011",
X=>mulr_2_91);

mulr_1_92<=a_1;
mulc_2_92 : entity work.gfmul
port map(
a=>a_2,
b=>"01011011",
X=>mulr_2_92);

mulr_1_93<=a_1;
mulc_2_93 : entity work.gfmul
port map(
a=>a_2,
b=>"10110110",
X=>mulr_2_93);

mulr_1_94<=a_1;
mulc_2_94 : entity work.gfmul
port map(
a=>a_2,
b=>"01110001",
X=>mulr_2_94);

mulr_1_95<=a_1;
mulc_2_95 : entity work.gfmul
port map(
a=>a_2,
b=>"11100010",
X=>mulr_2_95);

mulr_1_96<=a_1;
mulc_2_96 : entity work.gfmul
port map(
a=>a_2,
b=>"11011001",
X=>mulr_2_96);

mulr_1_97<=a_1;
mulc_2_97 : entity work.gfmul
port map(
a=>a_2,
b=>"10101111",
X=>mulr_2_97);

mulr_1_98<=a_1;
mulc_2_98 : entity work.gfmul
port map(
a=>a_2,
b=>"01000011",
X=>mulr_2_98);

mulr_1_99<=a_1;
mulc_2_99 : entity work.gfmul
port map(
a=>a_2,
b=>"10000110",
X=>mulr_2_99);

mulr_1_100<=a_1;
mulc_2_100 : entity work.gfmul
port map(
a=>a_2,
b=>"00010001",
X=>mulr_2_100);

mulr_1_101<=a_1;
mulc_2_101 : entity work.gfmul
port map(
a=>a_2,
b=>"00100010",
X=>mulr_2_101);

mulr_1_102<=a_1;
mulc_2_102 : entity work.gfmul
port map(
a=>a_2,
b=>"01000100",
X=>mulr_2_102);

mulr_1_103<=a_1;
mulc_2_103 : entity work.gfmul
port map(
a=>a_2,
b=>"10001000",
X=>mulr_2_103);

mulr_1_104<=a_1;
mulc_2_104 : entity work.gfmul
port map(
a=>a_2,
b=>"00001101",
X=>mulr_2_104);

mulr_1_105<=a_1;
mulc_2_105 : entity work.gfmul
port map(
a=>a_2,
b=>"00011010",
X=>mulr_2_105);

mulr_1_106<=a_1;
mulc_2_106 : entity work.gfmul
port map(
a=>a_2,
b=>"00110100",
X=>mulr_2_106);

mulr_1_107<=a_1;
mulc_2_107 : entity work.gfmul
port map(
a=>a_2,
b=>"01101000",
X=>mulr_2_107);

mulr_1_108<=a_1;
mulc_2_108 : entity work.gfmul
port map(
a=>a_2,
b=>"11010000",
X=>mulr_2_108);

mulr_1_109<=a_1;
mulc_2_109 : entity work.gfmul
port map(
a=>a_2,
b=>"10111101",
X=>mulr_2_109);

mulr_1_110<=a_1;
mulc_2_110 : entity work.gfmul
port map(
a=>a_2,
b=>"01100111",
X=>mulr_2_110);

mulr_1_111<=a_1;
mulc_2_111 : entity work.gfmul
port map(
a=>a_2,
b=>"11001110",
X=>mulr_2_111);

mulr_1_112<=a_1;
mulc_2_112 : entity work.gfmul
port map(
a=>a_2,
b=>"10000001",
X=>mulr_2_112);

mulr_1_113<=a_1;
mulc_2_113 : entity work.gfmul
port map(
a=>a_2,
b=>"00011111",
X=>mulr_2_113);

mulr_1_114<=a_1;
mulc_2_114 : entity work.gfmul
port map(
a=>a_2,
b=>"00111110",
X=>mulr_2_114);

mulr_1_115<=a_1;
mulc_2_115 : entity work.gfmul
port map(
a=>a_2,
b=>"01111100",
X=>mulr_2_115);

mulr_1_116<=a_1;
mulc_2_116 : entity work.gfmul
port map(
a=>a_2,
b=>"11111000",
X=>mulr_2_116);

mulr_1_117<=a_1;
mulc_2_117 : entity work.gfmul
port map(
a=>a_2,
b=>"11101101",
X=>mulr_2_117);

mulr_1_118<=a_1;
mulc_2_118 : entity work.gfmul
port map(
a=>a_2,
b=>"11000111",
X=>mulr_2_118);

mulr_1_119<=a_1;
mulc_2_119 : entity work.gfmul
port map(
a=>a_2,
b=>"10010011",
X=>mulr_2_119);

mulr_1_120<=a_1;
mulc_2_120 : entity work.gfmul
port map(
a=>a_2,
b=>"00111011",
X=>mulr_2_120);

mulr_1_121<=a_1;
mulc_2_121 : entity work.gfmul
port map(
a=>a_2,
b=>"01110110",
X=>mulr_2_121);

mulr_1_122<=a_1;
mulc_2_122 : entity work.gfmul
port map(
a=>a_2,
b=>"11101100",
X=>mulr_2_122);

mulr_1_123<=a_1;
mulc_2_123 : entity work.gfmul
port map(
a=>a_2,
b=>"11000101",
X=>mulr_2_123);

mulr_1_124<=a_1;
mulc_2_124 : entity work.gfmul
port map(
a=>a_2,
b=>"10010111",
X=>mulr_2_124);

mulr_1_125<=a_1;
mulc_2_125 : entity work.gfmul
port map(
a=>a_2,
b=>"00110011",
X=>mulr_2_125);

mulr_1_126<=a_1;
mulc_2_126 : entity work.gfmul
port map(
a=>a_2,
b=>"01100110",
X=>mulr_2_126);

mulr_1_127<=a_1;
mulc_2_127 : entity work.gfmul
port map(
a=>a_2,
b=>"11001100",
X=>mulr_2_127);

mulr_1_128<=a_1;
mulc_2_128 : entity work.gfmul
port map(
a=>a_2,
b=>"10000101",
X=>mulr_2_128);

mulr_1_129<=a_1;
mulc_2_129 : entity work.gfmul
port map(
a=>a_2,
b=>"00010111",
X=>mulr_2_129);

mulr_1_130<=a_1;
mulc_2_130 : entity work.gfmul
port map(
a=>a_2,
b=>"00101110",
X=>mulr_2_130);

mulr_1_131<=a_1;
mulc_2_131 : entity work.gfmul
port map(
a=>a_2,
b=>"01011100",
X=>mulr_2_131);

mulr_1_132<=a_1;
mulc_2_132 : entity work.gfmul
port map(
a=>a_2,
b=>"10111000",
X=>mulr_2_132);

mulr_1_133<=a_1;
mulc_2_133 : entity work.gfmul
port map(
a=>a_2,
b=>"01101101",
X=>mulr_2_133);

mulr_1_134<=a_1;
mulc_2_134 : entity work.gfmul
port map(
a=>a_2,
b=>"11011010",
X=>mulr_2_134);

mulr_1_135<=a_1;
mulc_2_135 : entity work.gfmul
port map(
a=>a_2,
b=>"10101001",
X=>mulr_2_135);

mulr_1_136<=a_1;
mulc_2_136 : entity work.gfmul
port map(
a=>a_2,
b=>"01001111",
X=>mulr_2_136);

mulr_1_137<=a_1;
mulc_2_137 : entity work.gfmul
port map(
a=>a_2,
b=>"10011110",
X=>mulr_2_137);

mulr_1_138<=a_1;
mulc_2_138 : entity work.gfmul
port map(
a=>a_2,
b=>"00100001",
X=>mulr_2_138);

mulr_1_139<=a_1;
mulc_2_139 : entity work.gfmul
port map(
a=>a_2,
b=>"01000010",
X=>mulr_2_139);

mulr_1_140<=a_1;
mulc_2_140 : entity work.gfmul
port map(
a=>a_2,
b=>"10000100",
X=>mulr_2_140);

mulr_1_141<=a_1;
mulc_2_141 : entity work.gfmul
port map(
a=>a_2,
b=>"00010101",
X=>mulr_2_141);

mulr_1_142<=a_1;
mulc_2_142 : entity work.gfmul
port map(
a=>a_2,
b=>"00101010",
X=>mulr_2_142);

mulr_1_143<=a_1;
mulc_2_143 : entity work.gfmul
port map(
a=>a_2,
b=>"01010100",
X=>mulr_2_143);

mulr_1_144<=a_1;
mulc_2_144 : entity work.gfmul
port map(
a=>a_2,
b=>"10101000",
X=>mulr_2_144);

mulr_1_145<=a_1;
mulc_2_145 : entity work.gfmul
port map(
a=>a_2,
b=>"01001101",
X=>mulr_2_145);

mulr_1_146<=a_1;
mulc_2_146 : entity work.gfmul
port map(
a=>a_2,
b=>"10011010",
X=>mulr_2_146);

mulr_1_147<=a_1;
mulc_2_147 : entity work.gfmul
port map(
a=>a_2,
b=>"00101001",
X=>mulr_2_147);

mulr_1_148<=a_1;
mulc_2_148 : entity work.gfmul
port map(
a=>a_2,
b=>"01010010",
X=>mulr_2_148);

mulr_1_149<=a_1;
mulc_2_149 : entity work.gfmul
port map(
a=>a_2,
b=>"10100100",
X=>mulr_2_149);

mulr_1_150<=a_1;
mulc_2_150 : entity work.gfmul
port map(
a=>a_2,
b=>"01010101",
X=>mulr_2_150);

mulr_1_151<=a_1;
mulc_2_151 : entity work.gfmul
port map(
a=>a_2,
b=>"10101010",
X=>mulr_2_151);

mulr_1_152<=a_1;
mulc_2_152 : entity work.gfmul
port map(
a=>a_2,
b=>"01001001",
X=>mulr_2_152);

mulr_1_153<=a_1;
mulc_2_153 : entity work.gfmul
port map(
a=>a_2,
b=>"10010010",
X=>mulr_2_153);

mulr_1_154<=a_1;
mulc_2_154 : entity work.gfmul
port map(
a=>a_2,
b=>"00111001",
X=>mulr_2_154);

mulr_1_155<=a_1;
mulc_2_155 : entity work.gfmul
port map(
a=>a_2,
b=>"01110010",
X=>mulr_2_155);

mulr_1_156<=a_1;
mulc_2_156 : entity work.gfmul
port map(
a=>a_2,
b=>"11100100",
X=>mulr_2_156);

mulr_1_157<=a_1;
mulc_2_157 : entity work.gfmul
port map(
a=>a_2,
b=>"11010101",
X=>mulr_2_157);

mulr_1_158<=a_1;
mulc_2_158 : entity work.gfmul
port map(
a=>a_2,
b=>"10110111",
X=>mulr_2_158);

mulr_1_159<=a_1;
mulc_2_159 : entity work.gfmul
port map(
a=>a_2,
b=>"01110011",
X=>mulr_2_159);

mulr_1_160<=a_1;
mulc_2_160 : entity work.gfmul
port map(
a=>a_2,
b=>"11100110",
X=>mulr_2_160);

mulr_1_161<=a_1;
mulc_2_161 : entity work.gfmul
port map(
a=>a_2,
b=>"11010001",
X=>mulr_2_161);

mulr_1_162<=a_1;
mulc_2_162 : entity work.gfmul
port map(
a=>a_2,
b=>"10111111",
X=>mulr_2_162);

mulr_1_163<=a_1;
mulc_2_163 : entity work.gfmul
port map(
a=>a_2,
b=>"01100011",
X=>mulr_2_163);

mulr_1_164<=a_1;
mulc_2_164 : entity work.gfmul
port map(
a=>a_2,
b=>"11000110",
X=>mulr_2_164);

mulr_1_165<=a_1;
mulc_2_165 : entity work.gfmul
port map(
a=>a_2,
b=>"10010001",
X=>mulr_2_165);

mulr_1_166<=a_1;
mulc_2_166 : entity work.gfmul
port map(
a=>a_2,
b=>"00111111",
X=>mulr_2_166);

mulr_1_167<=a_1;
mulc_2_167 : entity work.gfmul
port map(
a=>a_2,
b=>"01111110",
X=>mulr_2_167);

mulr_1_168<=a_1;
mulc_2_168 : entity work.gfmul
port map(
a=>a_2,
b=>"11111100",
X=>mulr_2_168);

mulr_1_169<=a_1;
mulc_2_169 : entity work.gfmul
port map(
a=>a_2,
b=>"11100101",
X=>mulr_2_169);

mulr_1_170<=a_1;
mulc_2_170 : entity work.gfmul
port map(
a=>a_2,
b=>"11010111",
X=>mulr_2_170);

mulr_1_171<=a_1;
mulc_2_171 : entity work.gfmul
port map(
a=>a_2,
b=>"10110011",
X=>mulr_2_171);

mulr_1_172<=a_1;
mulc_2_172 : entity work.gfmul
port map(
a=>a_2,
b=>"01111011",
X=>mulr_2_172);

mulr_1_173<=a_1;
mulc_2_173 : entity work.gfmul
port map(
a=>a_2,
b=>"11110110",
X=>mulr_2_173);

mulr_1_174<=a_1;
mulc_2_174 : entity work.gfmul
port map(
a=>a_2,
b=>"11110001",
X=>mulr_2_174);

mulr_1_175<=a_1;
mulc_2_175 : entity work.gfmul
port map(
a=>a_2,
b=>"11111111",
X=>mulr_2_175);

mulr_1_176<=a_1;
mulc_2_176 : entity work.gfmul
port map(
a=>a_2,
b=>"11100011",
X=>mulr_2_176);

mulr_1_177<=a_1;
mulc_2_177 : entity work.gfmul
port map(
a=>a_2,
b=>"11011011",
X=>mulr_2_177);

mulr_1_178<=a_1;
mulc_2_178 : entity work.gfmul
port map(
a=>a_2,
b=>"10101011",
X=>mulr_2_178);

mulr_1_179<=a_1;
mulc_2_179 : entity work.gfmul
port map(
a=>a_2,
b=>"01001011",
X=>mulr_2_179);

mulr_1_180<=a_1;
mulc_2_180 : entity work.gfmul
port map(
a=>a_2,
b=>"10010110",
X=>mulr_2_180);

mulr_1_181<=a_1;
mulc_2_181 : entity work.gfmul
port map(
a=>a_2,
b=>"00110001",
X=>mulr_2_181);

mulr_1_182<=a_1;
mulc_2_182 : entity work.gfmul
port map(
a=>a_2,
b=>"01100010",
X=>mulr_2_182);

mulr_1_183<=a_1;
mulc_2_183 : entity work.gfmul
port map(
a=>a_2,
b=>"11000100",
X=>mulr_2_183);

mulr_1_184<=a_1;
mulc_2_184 : entity work.gfmul
port map(
a=>a_2,
b=>"10010101",
X=>mulr_2_184);

mulr_1_185<=a_1;
mulc_2_185 : entity work.gfmul
port map(
a=>a_2,
b=>"00110111",
X=>mulr_2_185);

mulr_1_186<=a_1;
mulc_2_186 : entity work.gfmul
port map(
a=>a_2,
b=>"01101110",
X=>mulr_2_186);

mulr_1_187<=a_1;
mulc_2_187 : entity work.gfmul
port map(
a=>a_2,
b=>"11011100",
X=>mulr_2_187);

mulr_1_188<=a_1;
mulc_2_188 : entity work.gfmul
port map(
a=>a_2,
b=>"10100101",
X=>mulr_2_188);

mulr_1_189<=a_1;
mulc_2_189 : entity work.gfmul
port map(
a=>a_2,
b=>"01010111",
X=>mulr_2_189);

mulr_1_190<=a_1;
mulc_2_190 : entity work.gfmul
port map(
a=>a_2,
b=>"10101110",
X=>mulr_2_190);

mulr_1_191<=a_1;
mulc_2_191 : entity work.gfmul
port map(
a=>a_2,
b=>"01000001",
X=>mulr_2_191);

mulr_1_192<=a_1;
mulc_2_192 : entity work.gfmul
port map(
a=>a_2,
b=>"10000010",
X=>mulr_2_192);

mulr_1_193<=a_1;
mulc_2_193 : entity work.gfmul
port map(
a=>a_2,
b=>"00011001",
X=>mulr_2_193);

mulr_1_194<=a_1;
mulc_2_194 : entity work.gfmul
port map(
a=>a_2,
b=>"00110010",
X=>mulr_2_194);

mulr_1_195<=a_1;
mulc_2_195 : entity work.gfmul
port map(
a=>a_2,
b=>"01100100",
X=>mulr_2_195);

mulr_1_196<=a_1;
mulc_2_196 : entity work.gfmul
port map(
a=>a_2,
b=>"11001000",
X=>mulr_2_196);

mulr_1_197<=a_1;
mulc_2_197 : entity work.gfmul
port map(
a=>a_2,
b=>"10001101",
X=>mulr_2_197);

mulr_1_198<=a_1;
mulc_2_198 : entity work.gfmul
port map(
a=>a_2,
b=>"00000111",
X=>mulr_2_198);

mulr_1_199<=a_1;
mulc_2_199 : entity work.gfmul
port map(
a=>a_2,
b=>"00001110",
X=>mulr_2_199);

mulr_1_200<=a_1;
mulc_2_200 : entity work.gfmul
port map(
a=>a_2,
b=>"00011100",
X=>mulr_2_200);

mulr_1_201<=a_1;
mulc_2_201 : entity work.gfmul
port map(
a=>a_2,
b=>"00111000",
X=>mulr_2_201);

mulr_1_202<=a_1;
mulc_2_202 : entity work.gfmul
port map(
a=>a_2,
b=>"01110000",
X=>mulr_2_202);

mulr_1_203<=a_1;
mulc_2_203 : entity work.gfmul
port map(
a=>a_2,
b=>"11100000",
X=>mulr_2_203);

mulr_1_204<=a_1;
mulc_2_204 : entity work.gfmul
port map(
a=>a_2,
b=>"11011101",
X=>mulr_2_204);

mulr_1_205<=a_1;
mulc_2_205 : entity work.gfmul
port map(
a=>a_2,
b=>"10100111",
X=>mulr_2_205);

mulr_1_206<=a_1;
mulc_2_206 : entity work.gfmul
port map(
a=>a_2,
b=>"01010011",
X=>mulr_2_206);

mulr_1_207<=a_1;
mulc_2_207 : entity work.gfmul
port map(
a=>a_2,
b=>"10100110",
X=>mulr_2_207);

mulr_1_208<=a_1;
mulc_2_208 : entity work.gfmul
port map(
a=>a_2,
b=>"01010001",
X=>mulr_2_208);

mulr_1_209<=a_1;
mulc_2_209 : entity work.gfmul
port map(
a=>a_2,
b=>"10100010",
X=>mulr_2_209);

mulr_1_210<=a_1;
mulc_2_210 : entity work.gfmul
port map(
a=>a_2,
b=>"01011001",
X=>mulr_2_210);

mulr_1_211<=a_1;
mulc_2_211 : entity work.gfmul
port map(
a=>a_2,
b=>"10110010",
X=>mulr_2_211);

mulr_1_212<=a_1;
mulc_2_212 : entity work.gfmul
port map(
a=>a_2,
b=>"01111001",
X=>mulr_2_212);

mulr_1_213<=a_1;
mulc_2_213 : entity work.gfmul
port map(
a=>a_2,
b=>"11110010",
X=>mulr_2_213);

mulr_1_214<=a_1;
mulc_2_214 : entity work.gfmul
port map(
a=>a_2,
b=>"11111001",
X=>mulr_2_214);

mulr_1_215<=a_1;
mulc_2_215 : entity work.gfmul
port map(
a=>a_2,
b=>"11101111",
X=>mulr_2_215);

mulr_1_216<=a_1;
mulc_2_216 : entity work.gfmul
port map(
a=>a_2,
b=>"11000011",
X=>mulr_2_216);

mulr_1_217<=a_1;
mulc_2_217 : entity work.gfmul
port map(
a=>a_2,
b=>"10011011",
X=>mulr_2_217);

mulr_1_218<=a_1;
mulc_2_218 : entity work.gfmul
port map(
a=>a_2,
b=>"00101011",
X=>mulr_2_218);

mulr_1_219<=a_1;
mulc_2_219 : entity work.gfmul
port map(
a=>a_2,
b=>"01010110",
X=>mulr_2_219);

mulr_1_220<=a_1;
mulc_2_220 : entity work.gfmul
port map(
a=>a_2,
b=>"10101100",
X=>mulr_2_220);

mulr_1_221<=a_1;
mulc_2_221 : entity work.gfmul
port map(
a=>a_2,
b=>"01000101",
X=>mulr_2_221);

mulr_1_222<=a_1;
mulc_2_222 : entity work.gfmul
port map(
a=>a_2,
b=>"10001010",
X=>mulr_2_222);

mulr_1_223<=a_1;
mulc_2_223 : entity work.gfmul
port map(
a=>a_2,
b=>"00001001",
X=>mulr_2_223);

mulr_1_224<=a_1;
mulc_2_224 : entity work.gfmul
port map(
a=>a_2,
b=>"00010010",
X=>mulr_2_224);

mulr_1_225<=a_1;
mulc_2_225 : entity work.gfmul
port map(
a=>a_2,
b=>"00100100",
X=>mulr_2_225);

mulr_1_226<=a_1;
mulc_2_226 : entity work.gfmul
port map(
a=>a_2,
b=>"01001000",
X=>mulr_2_226);

mulr_1_227<=a_1;
mulc_2_227 : entity work.gfmul
port map(
a=>a_2,
b=>"10010000",
X=>mulr_2_227);

mulr_1_228<=a_1;
mulc_2_228 : entity work.gfmul
port map(
a=>a_2,
b=>"00111101",
X=>mulr_2_228);

mulr_1_229<=a_1;
mulc_2_229 : entity work.gfmul
port map(
a=>a_2,
b=>"01111010",
X=>mulr_2_229);

mulr_1_230<=a_1;
mulc_2_230 : entity work.gfmul
port map(
a=>a_2,
b=>"11110100",
X=>mulr_2_230);

mulr_1_231<=a_1;
mulc_2_231 : entity work.gfmul
port map(
a=>a_2,
b=>"11110101",
X=>mulr_2_231);

mulr_1_232<=a_1;
mulc_2_232 : entity work.gfmul
port map(
a=>a_2,
b=>"11110111",
X=>mulr_2_232);

mulr_1_233<=a_1;
mulc_2_233 : entity work.gfmul
port map(
a=>a_2,
b=>"11110011",
X=>mulr_2_233);

mulr_1_234<=a_1;
mulc_2_234 : entity work.gfmul
port map(
a=>a_2,
b=>"11111011",
X=>mulr_2_234);

mulr_1_235<=a_1;
mulc_2_235 : entity work.gfmul
port map(
a=>a_2,
b=>"11101011",
X=>mulr_2_235);

mulr_1_236<=a_1;
mulc_2_236 : entity work.gfmul
port map(
a=>a_2,
b=>"11001011",
X=>mulr_2_236);

mulr_1_237<=a_1;
mulc_2_237 : entity work.gfmul
port map(
a=>a_2,
b=>"10001011",
X=>mulr_2_237);

mulr_1_238<=a_1;
mulc_2_238 : entity work.gfmul
port map(
a=>a_2,
b=>"00001011",
X=>mulr_2_238);

mulr_1_239<=a_1;
mulc_2_239 : entity work.gfmul
port map(
a=>a_2,
b=>"00010110",
X=>mulr_2_239);

mulr_1_240<=a_1;
mulc_2_240 : entity work.gfmul
port map(
a=>a_2,
b=>"00101100",
X=>mulr_2_240);

mulr_1_241<=a_1;
mulc_2_241 : entity work.gfmul
port map(
a=>a_2,
b=>"01011000",
X=>mulr_2_241);

mulr_1_242<=a_1;
mulc_2_242 : entity work.gfmul
port map(
a=>a_2,
b=>"10110000",
X=>mulr_2_242);

mulr_1_243<=a_1;
mulc_2_243 : entity work.gfmul
port map(
a=>a_2,
b=>"01111101",
X=>mulr_2_243);

mulr_1_244<=a_1;
mulc_2_244 : entity work.gfmul
port map(
a=>a_2,
b=>"11111010",
X=>mulr_2_244);

mulr_1_245<=a_1;
mulc_2_245 : entity work.gfmul
port map(
a=>a_2,
b=>"11101001",
X=>mulr_2_245);

mulr_1_246<=a_1;
mulc_2_246 : entity work.gfmul
port map(
a=>a_2,
b=>"11001111",
X=>mulr_2_246);

mulr_1_247<=a_1;
mulc_2_247 : entity work.gfmul
port map(
a=>a_2,
b=>"10000011",
X=>mulr_2_247);

mulr_1_248<=a_1;
mulc_2_248 : entity work.gfmul
port map(
a=>a_2,
b=>"00011011",
X=>mulr_2_248);

mulr_1_249<=a_1;
mulc_2_249 : entity work.gfmul
port map(
a=>a_2,
b=>"00110110",
X=>mulr_2_249);

mulr_1_250<=a_1;
mulc_2_250 : entity work.gfmul
port map(
a=>a_2,
b=>"01101100",
X=>mulr_2_250);

mulr_1_251<=a_1;
mulc_2_251 : entity work.gfmul
port map(
a=>a_2,
b=>"11011000",
X=>mulr_2_251);

mulr_1_252<=a_1;
mulc_2_252 : entity work.gfmul
port map(
a=>a_2,
b=>"10101101",
X=>mulr_2_252);

mulr_1_253<=a_1;
mulc_2_253 : entity work.gfmul
port map(
a=>a_2,
b=>"01000111",
X=>mulr_2_253);

mulr_1_254<=a_1;
mulc_2_254 : entity work.gfmul
port map(
a=>a_2,
b=>"10001110",
X=>mulr_2_254);

mulr_1_255<=a_1;
mulc_2_255 : entity work.gfmul
port map(
a=>a_2,
b=>"00000001",
X=>mulr_2_255);

sumr_1<= mulr_1_1 xor mulr_2_1;
sumr_2<= mulr_1_2 xor mulr_2_2;
sumr_3<= mulr_1_3 xor mulr_2_3;
sumr_4<= mulr_1_4 xor mulr_2_4;
sumr_5<= mulr_1_5 xor mulr_2_5;
sumr_6<= mulr_1_6 xor mulr_2_6;
sumr_7<= mulr_1_7 xor mulr_2_7;
sumr_8<= mulr_1_8 xor mulr_2_8;
sumr_9<= mulr_1_9 xor mulr_2_9;
sumr_10<= mulr_1_10 xor mulr_2_10;
sumr_11<= mulr_1_11 xor mulr_2_11;
sumr_12<= mulr_1_12 xor mulr_2_12;
sumr_13<= mulr_1_13 xor mulr_2_13;
sumr_14<= mulr_1_14 xor mulr_2_14;
sumr_15<= mulr_1_15 xor mulr_2_15;
sumr_16<= mulr_1_16 xor mulr_2_16;
sumr_17<= mulr_1_17 xor mulr_2_17;
sumr_18<= mulr_1_18 xor mulr_2_18;
sumr_19<= mulr_1_19 xor mulr_2_19;
sumr_20<= mulr_1_20 xor mulr_2_20;
sumr_21<= mulr_1_21 xor mulr_2_21;
sumr_22<= mulr_1_22 xor mulr_2_22;
sumr_23<= mulr_1_23 xor mulr_2_23;
sumr_24<= mulr_1_24 xor mulr_2_24;
sumr_25<= mulr_1_25 xor mulr_2_25;
sumr_26<= mulr_1_26 xor mulr_2_26;
sumr_27<= mulr_1_27 xor mulr_2_27;
sumr_28<= mulr_1_28 xor mulr_2_28;
sumr_29<= mulr_1_29 xor mulr_2_29;
sumr_30<= mulr_1_30 xor mulr_2_30;
sumr_31<= mulr_1_31 xor mulr_2_31;
sumr_32<= mulr_1_32 xor mulr_2_32;
sumr_33<= mulr_1_33 xor mulr_2_33;
sumr_34<= mulr_1_34 xor mulr_2_34;
sumr_35<= mulr_1_35 xor mulr_2_35;
sumr_36<= mulr_1_36 xor mulr_2_36;
sumr_37<= mulr_1_37 xor mulr_2_37;
sumr_38<= mulr_1_38 xor mulr_2_38;
sumr_39<= mulr_1_39 xor mulr_2_39;
sumr_40<= mulr_1_40 xor mulr_2_40;
sumr_41<= mulr_1_41 xor mulr_2_41;
sumr_42<= mulr_1_42 xor mulr_2_42;
sumr_43<= mulr_1_43 xor mulr_2_43;
sumr_44<= mulr_1_44 xor mulr_2_44;
sumr_45<= mulr_1_45 xor mulr_2_45;
sumr_46<= mulr_1_46 xor mulr_2_46;
sumr_47<= mulr_1_47 xor mulr_2_47;
sumr_48<= mulr_1_48 xor mulr_2_48;
sumr_49<= mulr_1_49 xor mulr_2_49;
sumr_50<= mulr_1_50 xor mulr_2_50;
sumr_51<= mulr_1_51 xor mulr_2_51;
sumr_52<= mulr_1_52 xor mulr_2_52;
sumr_53<= mulr_1_53 xor mulr_2_53;
sumr_54<= mulr_1_54 xor mulr_2_54;
sumr_55<= mulr_1_55 xor mulr_2_55;
sumr_56<= mulr_1_56 xor mulr_2_56;
sumr_57<= mulr_1_57 xor mulr_2_57;
sumr_58<= mulr_1_58 xor mulr_2_58;
sumr_59<= mulr_1_59 xor mulr_2_59;
sumr_60<= mulr_1_60 xor mulr_2_60;
sumr_61<= mulr_1_61 xor mulr_2_61;
sumr_62<= mulr_1_62 xor mulr_2_62;
sumr_63<= mulr_1_63 xor mulr_2_63;
sumr_64<= mulr_1_64 xor mulr_2_64;
sumr_65<= mulr_1_65 xor mulr_2_65;
sumr_66<= mulr_1_66 xor mulr_2_66;
sumr_67<= mulr_1_67 xor mulr_2_67;
sumr_68<= mulr_1_68 xor mulr_2_68;
sumr_69<= mulr_1_69 xor mulr_2_69;
sumr_70<= mulr_1_70 xor mulr_2_70;
sumr_71<= mulr_1_71 xor mulr_2_71;
sumr_72<= mulr_1_72 xor mulr_2_72;
sumr_73<= mulr_1_73 xor mulr_2_73;
sumr_74<= mulr_1_74 xor mulr_2_74;
sumr_75<= mulr_1_75 xor mulr_2_75;
sumr_76<= mulr_1_76 xor mulr_2_76;
sumr_77<= mulr_1_77 xor mulr_2_77;
sumr_78<= mulr_1_78 xor mulr_2_78;
sumr_79<= mulr_1_79 xor mulr_2_79;
sumr_80<= mulr_1_80 xor mulr_2_80;
sumr_81<= mulr_1_81 xor mulr_2_81;
sumr_82<= mulr_1_82 xor mulr_2_82;
sumr_83<= mulr_1_83 xor mulr_2_83;
sumr_84<= mulr_1_84 xor mulr_2_84;
sumr_85<= mulr_1_85 xor mulr_2_85;
sumr_86<= mulr_1_86 xor mulr_2_86;
sumr_87<= mulr_1_87 xor mulr_2_87;
sumr_88<= mulr_1_88 xor mulr_2_88;
sumr_89<= mulr_1_89 xor mulr_2_89;
sumr_90<= mulr_1_90 xor mulr_2_90;
sumr_91<= mulr_1_91 xor mulr_2_91;
sumr_92<= mulr_1_92 xor mulr_2_92;
sumr_93<= mulr_1_93 xor mulr_2_93;
sumr_94<= mulr_1_94 xor mulr_2_94;
sumr_95<= mulr_1_95 xor mulr_2_95;
sumr_96<= mulr_1_96 xor mulr_2_96;
sumr_97<= mulr_1_97 xor mulr_2_97;
sumr_98<= mulr_1_98 xor mulr_2_98;
sumr_99<= mulr_1_99 xor mulr_2_99;
sumr_100<= mulr_1_100 xor mulr_2_100;
sumr_101<= mulr_1_101 xor mulr_2_101;
sumr_102<= mulr_1_102 xor mulr_2_102;
sumr_103<= mulr_1_103 xor mulr_2_103;
sumr_104<= mulr_1_104 xor mulr_2_104;
sumr_105<= mulr_1_105 xor mulr_2_105;
sumr_106<= mulr_1_106 xor mulr_2_106;
sumr_107<= mulr_1_107 xor mulr_2_107;
sumr_108<= mulr_1_108 xor mulr_2_108;
sumr_109<= mulr_1_109 xor mulr_2_109;
sumr_110<= mulr_1_110 xor mulr_2_110;
sumr_111<= mulr_1_111 xor mulr_2_111;
sumr_112<= mulr_1_112 xor mulr_2_112;
sumr_113<= mulr_1_113 xor mulr_2_113;
sumr_114<= mulr_1_114 xor mulr_2_114;
sumr_115<= mulr_1_115 xor mulr_2_115;
sumr_116<= mulr_1_116 xor mulr_2_116;
sumr_117<= mulr_1_117 xor mulr_2_117;
sumr_118<= mulr_1_118 xor mulr_2_118;
sumr_119<= mulr_1_119 xor mulr_2_119;
sumr_120<= mulr_1_120 xor mulr_2_120;
sumr_121<= mulr_1_121 xor mulr_2_121;
sumr_122<= mulr_1_122 xor mulr_2_122;
sumr_123<= mulr_1_123 xor mulr_2_123;
sumr_124<= mulr_1_124 xor mulr_2_124;
sumr_125<= mulr_1_125 xor mulr_2_125;
sumr_126<= mulr_1_126 xor mulr_2_126;
sumr_127<= mulr_1_127 xor mulr_2_127;
sumr_128<= mulr_1_128 xor mulr_2_128;
sumr_129<= mulr_1_129 xor mulr_2_129;
sumr_130<= mulr_1_130 xor mulr_2_130;
sumr_131<= mulr_1_131 xor mulr_2_131;
sumr_132<= mulr_1_132 xor mulr_2_132;
sumr_133<= mulr_1_133 xor mulr_2_133;
sumr_134<= mulr_1_134 xor mulr_2_134;
sumr_135<= mulr_1_135 xor mulr_2_135;
sumr_136<= mulr_1_136 xor mulr_2_136;
sumr_137<= mulr_1_137 xor mulr_2_137;
sumr_138<= mulr_1_138 xor mulr_2_138;
sumr_139<= mulr_1_139 xor mulr_2_139;
sumr_140<= mulr_1_140 xor mulr_2_140;
sumr_141<= mulr_1_141 xor mulr_2_141;
sumr_142<= mulr_1_142 xor mulr_2_142;
sumr_143<= mulr_1_143 xor mulr_2_143;
sumr_144<= mulr_1_144 xor mulr_2_144;
sumr_145<= mulr_1_145 xor mulr_2_145;
sumr_146<= mulr_1_146 xor mulr_2_146;
sumr_147<= mulr_1_147 xor mulr_2_147;
sumr_148<= mulr_1_148 xor mulr_2_148;
sumr_149<= mulr_1_149 xor mulr_2_149;
sumr_150<= mulr_1_150 xor mulr_2_150;
sumr_151<= mulr_1_151 xor mulr_2_151;
sumr_152<= mulr_1_152 xor mulr_2_152;
sumr_153<= mulr_1_153 xor mulr_2_153;
sumr_154<= mulr_1_154 xor mulr_2_154;
sumr_155<= mulr_1_155 xor mulr_2_155;
sumr_156<= mulr_1_156 xor mulr_2_156;
sumr_157<= mulr_1_157 xor mulr_2_157;
sumr_158<= mulr_1_158 xor mulr_2_158;
sumr_159<= mulr_1_159 xor mulr_2_159;
sumr_160<= mulr_1_160 xor mulr_2_160;
sumr_161<= mulr_1_161 xor mulr_2_161;
sumr_162<= mulr_1_162 xor mulr_2_162;
sumr_163<= mulr_1_163 xor mulr_2_163;
sumr_164<= mulr_1_164 xor mulr_2_164;
sumr_165<= mulr_1_165 xor mulr_2_165;
sumr_166<= mulr_1_166 xor mulr_2_166;
sumr_167<= mulr_1_167 xor mulr_2_167;
sumr_168<= mulr_1_168 xor mulr_2_168;
sumr_169<= mulr_1_169 xor mulr_2_169;
sumr_170<= mulr_1_170 xor mulr_2_170;
sumr_171<= mulr_1_171 xor mulr_2_171;
sumr_172<= mulr_1_172 xor mulr_2_172;
sumr_173<= mulr_1_173 xor mulr_2_173;
sumr_174<= mulr_1_174 xor mulr_2_174;
sumr_175<= mulr_1_175 xor mulr_2_175;
sumr_176<= mulr_1_176 xor mulr_2_176;
sumr_177<= mulr_1_177 xor mulr_2_177;
sumr_178<= mulr_1_178 xor mulr_2_178;
sumr_179<= mulr_1_179 xor mulr_2_179;
sumr_180<= mulr_1_180 xor mulr_2_180;
sumr_181<= mulr_1_181 xor mulr_2_181;
sumr_182<= mulr_1_182 xor mulr_2_182;
sumr_183<= mulr_1_183 xor mulr_2_183;
sumr_184<= mulr_1_184 xor mulr_2_184;
sumr_185<= mulr_1_185 xor mulr_2_185;
sumr_186<= mulr_1_186 xor mulr_2_186;
sumr_187<= mulr_1_187 xor mulr_2_187;
sumr_188<= mulr_1_188 xor mulr_2_188;
sumr_189<= mulr_1_189 xor mulr_2_189;
sumr_190<= mulr_1_190 xor mulr_2_190;
sumr_191<= mulr_1_191 xor mulr_2_191;
sumr_192<= mulr_1_192 xor mulr_2_192;
sumr_193<= mulr_1_193 xor mulr_2_193;
sumr_194<= mulr_1_194 xor mulr_2_194;
sumr_195<= mulr_1_195 xor mulr_2_195;
sumr_196<= mulr_1_196 xor mulr_2_196;
sumr_197<= mulr_1_197 xor mulr_2_197;
sumr_198<= mulr_1_198 xor mulr_2_198;
sumr_199<= mulr_1_199 xor mulr_2_199;
sumr_200<= mulr_1_200 xor mulr_2_200;
sumr_201<= mulr_1_201 xor mulr_2_201;
sumr_202<= mulr_1_202 xor mulr_2_202;
sumr_203<= mulr_1_203 xor mulr_2_203;
sumr_204<= mulr_1_204 xor mulr_2_204;
sumr_205<= mulr_1_205 xor mulr_2_205;
sumr_206<= mulr_1_206 xor mulr_2_206;
sumr_207<= mulr_1_207 xor mulr_2_207;
sumr_208<= mulr_1_208 xor mulr_2_208;
sumr_209<= mulr_1_209 xor mulr_2_209;
sumr_210<= mulr_1_210 xor mulr_2_210;
sumr_211<= mulr_1_211 xor mulr_2_211;
sumr_212<= mulr_1_212 xor mulr_2_212;
sumr_213<= mulr_1_213 xor mulr_2_213;
sumr_214<= mulr_1_214 xor mulr_2_214;
sumr_215<= mulr_1_215 xor mulr_2_215;
sumr_216<= mulr_1_216 xor mulr_2_216;
sumr_217<= mulr_1_217 xor mulr_2_217;
sumr_218<= mulr_1_218 xor mulr_2_218;
sumr_219<= mulr_1_219 xor mulr_2_219;
sumr_220<= mulr_1_220 xor mulr_2_220;
sumr_221<= mulr_1_221 xor mulr_2_221;
sumr_222<= mulr_1_222 xor mulr_2_222;
sumr_223<= mulr_1_223 xor mulr_2_223;
sumr_224<= mulr_1_224 xor mulr_2_224;
sumr_225<= mulr_1_225 xor mulr_2_225;
sumr_226<= mulr_1_226 xor mulr_2_226;
sumr_227<= mulr_1_227 xor mulr_2_227;
sumr_228<= mulr_1_228 xor mulr_2_228;
sumr_229<= mulr_1_229 xor mulr_2_229;
sumr_230<= mulr_1_230 xor mulr_2_230;
sumr_231<= mulr_1_231 xor mulr_2_231;
sumr_232<= mulr_1_232 xor mulr_2_232;
sumr_233<= mulr_1_233 xor mulr_2_233;
sumr_234<= mulr_1_234 xor mulr_2_234;
sumr_235<= mulr_1_235 xor mulr_2_235;
sumr_236<= mulr_1_236 xor mulr_2_236;
sumr_237<= mulr_1_237 xor mulr_2_237;
sumr_238<= mulr_1_238 xor mulr_2_238;
sumr_239<= mulr_1_239 xor mulr_2_239;
sumr_240<= mulr_1_240 xor mulr_2_240;
sumr_241<= mulr_1_241 xor mulr_2_241;
sumr_242<= mulr_1_242 xor mulr_2_242;
sumr_243<= mulr_1_243 xor mulr_2_243;
sumr_244<= mulr_1_244 xor mulr_2_244;
sumr_245<= mulr_1_245 xor mulr_2_245;
sumr_246<= mulr_1_246 xor mulr_2_246;
sumr_247<= mulr_1_247 xor mulr_2_247;
sumr_248<= mulr_1_248 xor mulr_2_248;
sumr_249<= mulr_1_249 xor mulr_2_249;
sumr_250<= mulr_1_250 xor mulr_2_250;
sumr_251<= mulr_1_251 xor mulr_2_251;
sumr_252<= mulr_1_252 xor mulr_2_252;
sumr_253<= mulr_1_253 xor mulr_2_253;
sumr_254<= mulr_1_254 xor mulr_2_254;
sumr_255<= mulr_1_255 xor mulr_2_255;
E(254)<=not ( sumr_1(0) or sumr_1(1) or sumr_1(2) or sumr_1(3) or sumr_1(4) or sumr_1(5) or sumr_1(6) or sumr_1(7));
E(253)<=not ( sumr_2(0) or sumr_2(1) or sumr_2(2) or sumr_2(3) or sumr_2(4) or sumr_2(5) or sumr_2(6) or sumr_2(7));
E(252)<=not ( sumr_3(0) or sumr_3(1) or sumr_3(2) or sumr_3(3) or sumr_3(4) or sumr_3(5) or sumr_3(6) or sumr_3(7));
E(251)<=not ( sumr_4(0) or sumr_4(1) or sumr_4(2) or sumr_4(3) or sumr_4(4) or sumr_4(5) or sumr_4(6) or sumr_4(7));
E(250)<=not ( sumr_5(0) or sumr_5(1) or sumr_5(2) or sumr_5(3) or sumr_5(4) or sumr_5(5) or sumr_5(6) or sumr_5(7));
E(249)<=not ( sumr_6(0) or sumr_6(1) or sumr_6(2) or sumr_6(3) or sumr_6(4) or sumr_6(5) or sumr_6(6) or sumr_6(7));
E(248)<=not ( sumr_7(0) or sumr_7(1) or sumr_7(2) or sumr_7(3) or sumr_7(4) or sumr_7(5) or sumr_7(6) or sumr_7(7));
E(247)<=not ( sumr_8(0) or sumr_8(1) or sumr_8(2) or sumr_8(3) or sumr_8(4) or sumr_8(5) or sumr_8(6) or sumr_8(7));
E(246)<=not ( sumr_9(0) or sumr_9(1) or sumr_9(2) or sumr_9(3) or sumr_9(4) or sumr_9(5) or sumr_9(6) or sumr_9(7));
E(245)<=not ( sumr_10(0) or sumr_10(1) or sumr_10(2) or sumr_10(3) or sumr_10(4) or sumr_10(5) or sumr_10(6) or sumr_10(7));
E(244)<=not ( sumr_11(0) or sumr_11(1) or sumr_11(2) or sumr_11(3) or sumr_11(4) or sumr_11(5) or sumr_11(6) or sumr_11(7));
E(243)<=not ( sumr_12(0) or sumr_12(1) or sumr_12(2) or sumr_12(3) or sumr_12(4) or sumr_12(5) or sumr_12(6) or sumr_12(7));
E(242)<=not ( sumr_13(0) or sumr_13(1) or sumr_13(2) or sumr_13(3) or sumr_13(4) or sumr_13(5) or sumr_13(6) or sumr_13(7));
E(241)<=not ( sumr_14(0) or sumr_14(1) or sumr_14(2) or sumr_14(3) or sumr_14(4) or sumr_14(5) or sumr_14(6) or sumr_14(7));
E(240)<=not ( sumr_15(0) or sumr_15(1) or sumr_15(2) or sumr_15(3) or sumr_15(4) or sumr_15(5) or sumr_15(6) or sumr_15(7));
E(239)<=not ( sumr_16(0) or sumr_16(1) or sumr_16(2) or sumr_16(3) or sumr_16(4) or sumr_16(5) or sumr_16(6) or sumr_16(7));
E(238)<=not ( sumr_17(0) or sumr_17(1) or sumr_17(2) or sumr_17(3) or sumr_17(4) or sumr_17(5) or sumr_17(6) or sumr_17(7));
E(237)<=not ( sumr_18(0) or sumr_18(1) or sumr_18(2) or sumr_18(3) or sumr_18(4) or sumr_18(5) or sumr_18(6) or sumr_18(7));
E(236)<=not ( sumr_19(0) or sumr_19(1) or sumr_19(2) or sumr_19(3) or sumr_19(4) or sumr_19(5) or sumr_19(6) or sumr_19(7));
E(235)<=not ( sumr_20(0) or sumr_20(1) or sumr_20(2) or sumr_20(3) or sumr_20(4) or sumr_20(5) or sumr_20(6) or sumr_20(7));
E(234)<=not ( sumr_21(0) or sumr_21(1) or sumr_21(2) or sumr_21(3) or sumr_21(4) or sumr_21(5) or sumr_21(6) or sumr_21(7));
E(233)<=not ( sumr_22(0) or sumr_22(1) or sumr_22(2) or sumr_22(3) or sumr_22(4) or sumr_22(5) or sumr_22(6) or sumr_22(7));
E(232)<=not ( sumr_23(0) or sumr_23(1) or sumr_23(2) or sumr_23(3) or sumr_23(4) or sumr_23(5) or sumr_23(6) or sumr_23(7));
E(231)<=not ( sumr_24(0) or sumr_24(1) or sumr_24(2) or sumr_24(3) or sumr_24(4) or sumr_24(5) or sumr_24(6) or sumr_24(7));
E(230)<=not ( sumr_25(0) or sumr_25(1) or sumr_25(2) or sumr_25(3) or sumr_25(4) or sumr_25(5) or sumr_25(6) or sumr_25(7));
E(229)<=not ( sumr_26(0) or sumr_26(1) or sumr_26(2) or sumr_26(3) or sumr_26(4) or sumr_26(5) or sumr_26(6) or sumr_26(7));
E(228)<=not ( sumr_27(0) or sumr_27(1) or sumr_27(2) or sumr_27(3) or sumr_27(4) or sumr_27(5) or sumr_27(6) or sumr_27(7));
E(227)<=not ( sumr_28(0) or sumr_28(1) or sumr_28(2) or sumr_28(3) or sumr_28(4) or sumr_28(5) or sumr_28(6) or sumr_28(7));
E(226)<=not ( sumr_29(0) or sumr_29(1) or sumr_29(2) or sumr_29(3) or sumr_29(4) or sumr_29(5) or sumr_29(6) or sumr_29(7));
E(225)<=not ( sumr_30(0) or sumr_30(1) or sumr_30(2) or sumr_30(3) or sumr_30(4) or sumr_30(5) or sumr_30(6) or sumr_30(7));
E(224)<=not ( sumr_31(0) or sumr_31(1) or sumr_31(2) or sumr_31(3) or sumr_31(4) or sumr_31(5) or sumr_31(6) or sumr_31(7));
E(223)<=not ( sumr_32(0) or sumr_32(1) or sumr_32(2) or sumr_32(3) or sumr_32(4) or sumr_32(5) or sumr_32(6) or sumr_32(7));
E(222)<=not ( sumr_33(0) or sumr_33(1) or sumr_33(2) or sumr_33(3) or sumr_33(4) or sumr_33(5) or sumr_33(6) or sumr_33(7));
E(221)<=not ( sumr_34(0) or sumr_34(1) or sumr_34(2) or sumr_34(3) or sumr_34(4) or sumr_34(5) or sumr_34(6) or sumr_34(7));
E(220)<=not ( sumr_35(0) or sumr_35(1) or sumr_35(2) or sumr_35(3) or sumr_35(4) or sumr_35(5) or sumr_35(6) or sumr_35(7));
E(219)<=not ( sumr_36(0) or sumr_36(1) or sumr_36(2) or sumr_36(3) or sumr_36(4) or sumr_36(5) or sumr_36(6) or sumr_36(7));
E(218)<=not ( sumr_37(0) or sumr_37(1) or sumr_37(2) or sumr_37(3) or sumr_37(4) or sumr_37(5) or sumr_37(6) or sumr_37(7));
E(217)<=not ( sumr_38(0) or sumr_38(1) or sumr_38(2) or sumr_38(3) or sumr_38(4) or sumr_38(5) or sumr_38(6) or sumr_38(7));
E(216)<=not ( sumr_39(0) or sumr_39(1) or sumr_39(2) or sumr_39(3) or sumr_39(4) or sumr_39(5) or sumr_39(6) or sumr_39(7));
E(215)<=not ( sumr_40(0) or sumr_40(1) or sumr_40(2) or sumr_40(3) or sumr_40(4) or sumr_40(5) or sumr_40(6) or sumr_40(7));
E(214)<=not ( sumr_41(0) or sumr_41(1) or sumr_41(2) or sumr_41(3) or sumr_41(4) or sumr_41(5) or sumr_41(6) or sumr_41(7));
E(213)<=not ( sumr_42(0) or sumr_42(1) or sumr_42(2) or sumr_42(3) or sumr_42(4) or sumr_42(5) or sumr_42(6) or sumr_42(7));
E(212)<=not ( sumr_43(0) or sumr_43(1) or sumr_43(2) or sumr_43(3) or sumr_43(4) or sumr_43(5) or sumr_43(6) or sumr_43(7));
E(211)<=not ( sumr_44(0) or sumr_44(1) or sumr_44(2) or sumr_44(3) or sumr_44(4) or sumr_44(5) or sumr_44(6) or sumr_44(7));
E(210)<=not ( sumr_45(0) or sumr_45(1) or sumr_45(2) or sumr_45(3) or sumr_45(4) or sumr_45(5) or sumr_45(6) or sumr_45(7));
E(209)<=not ( sumr_46(0) or sumr_46(1) or sumr_46(2) or sumr_46(3) or sumr_46(4) or sumr_46(5) or sumr_46(6) or sumr_46(7));
E(208)<=not ( sumr_47(0) or sumr_47(1) or sumr_47(2) or sumr_47(3) or sumr_47(4) or sumr_47(5) or sumr_47(6) or sumr_47(7));
E(207)<=not ( sumr_48(0) or sumr_48(1) or sumr_48(2) or sumr_48(3) or sumr_48(4) or sumr_48(5) or sumr_48(6) or sumr_48(7));
E(206)<=not ( sumr_49(0) or sumr_49(1) or sumr_49(2) or sumr_49(3) or sumr_49(4) or sumr_49(5) or sumr_49(6) or sumr_49(7));
E(205)<=not ( sumr_50(0) or sumr_50(1) or sumr_50(2) or sumr_50(3) or sumr_50(4) or sumr_50(5) or sumr_50(6) or sumr_50(7));
E(204)<=not ( sumr_51(0) or sumr_51(1) or sumr_51(2) or sumr_51(3) or sumr_51(4) or sumr_51(5) or sumr_51(6) or sumr_51(7));
E(203)<=not ( sumr_52(0) or sumr_52(1) or sumr_52(2) or sumr_52(3) or sumr_52(4) or sumr_52(5) or sumr_52(6) or sumr_52(7));
E(202)<=not ( sumr_53(0) or sumr_53(1) or sumr_53(2) or sumr_53(3) or sumr_53(4) or sumr_53(5) or sumr_53(6) or sumr_53(7));
E(201)<=not ( sumr_54(0) or sumr_54(1) or sumr_54(2) or sumr_54(3) or sumr_54(4) or sumr_54(5) or sumr_54(6) or sumr_54(7));
E(200)<=not ( sumr_55(0) or sumr_55(1) or sumr_55(2) or sumr_55(3) or sumr_55(4) or sumr_55(5) or sumr_55(6) or sumr_55(7));
E(199)<=not ( sumr_56(0) or sumr_56(1) or sumr_56(2) or sumr_56(3) or sumr_56(4) or sumr_56(5) or sumr_56(6) or sumr_56(7));
E(198)<=not ( sumr_57(0) or sumr_57(1) or sumr_57(2) or sumr_57(3) or sumr_57(4) or sumr_57(5) or sumr_57(6) or sumr_57(7));
E(197)<=not ( sumr_58(0) or sumr_58(1) or sumr_58(2) or sumr_58(3) or sumr_58(4) or sumr_58(5) or sumr_58(6) or sumr_58(7));
E(196)<=not ( sumr_59(0) or sumr_59(1) or sumr_59(2) or sumr_59(3) or sumr_59(4) or sumr_59(5) or sumr_59(6) or sumr_59(7));
E(195)<=not ( sumr_60(0) or sumr_60(1) or sumr_60(2) or sumr_60(3) or sumr_60(4) or sumr_60(5) or sumr_60(6) or sumr_60(7));
E(194)<=not ( sumr_61(0) or sumr_61(1) or sumr_61(2) or sumr_61(3) or sumr_61(4) or sumr_61(5) or sumr_61(6) or sumr_61(7));
E(193)<=not ( sumr_62(0) or sumr_62(1) or sumr_62(2) or sumr_62(3) or sumr_62(4) or sumr_62(5) or sumr_62(6) or sumr_62(7));
E(192)<=not ( sumr_63(0) or sumr_63(1) or sumr_63(2) or sumr_63(3) or sumr_63(4) or sumr_63(5) or sumr_63(6) or sumr_63(7));
E(191)<=not ( sumr_64(0) or sumr_64(1) or sumr_64(2) or sumr_64(3) or sumr_64(4) or sumr_64(5) or sumr_64(6) or sumr_64(7));
E(190)<=not ( sumr_65(0) or sumr_65(1) or sumr_65(2) or sumr_65(3) or sumr_65(4) or sumr_65(5) or sumr_65(6) or sumr_65(7));
E(189)<=not ( sumr_66(0) or sumr_66(1) or sumr_66(2) or sumr_66(3) or sumr_66(4) or sumr_66(5) or sumr_66(6) or sumr_66(7));
E(188)<=not ( sumr_67(0) or sumr_67(1) or sumr_67(2) or sumr_67(3) or sumr_67(4) or sumr_67(5) or sumr_67(6) or sumr_67(7));
E(187)<=not ( sumr_68(0) or sumr_68(1) or sumr_68(2) or sumr_68(3) or sumr_68(4) or sumr_68(5) or sumr_68(6) or sumr_68(7));
E(186)<=not ( sumr_69(0) or sumr_69(1) or sumr_69(2) or sumr_69(3) or sumr_69(4) or sumr_69(5) or sumr_69(6) or sumr_69(7));
E(185)<=not ( sumr_70(0) or sumr_70(1) or sumr_70(2) or sumr_70(3) or sumr_70(4) or sumr_70(5) or sumr_70(6) or sumr_70(7));
E(184)<=not ( sumr_71(0) or sumr_71(1) or sumr_71(2) or sumr_71(3) or sumr_71(4) or sumr_71(5) or sumr_71(6) or sumr_71(7));
E(183)<=not ( sumr_72(0) or sumr_72(1) or sumr_72(2) or sumr_72(3) or sumr_72(4) or sumr_72(5) or sumr_72(6) or sumr_72(7));
E(182)<=not ( sumr_73(0) or sumr_73(1) or sumr_73(2) or sumr_73(3) or sumr_73(4) or sumr_73(5) or sumr_73(6) or sumr_73(7));
E(181)<=not ( sumr_74(0) or sumr_74(1) or sumr_74(2) or sumr_74(3) or sumr_74(4) or sumr_74(5) or sumr_74(6) or sumr_74(7));
E(180)<=not ( sumr_75(0) or sumr_75(1) or sumr_75(2) or sumr_75(3) or sumr_75(4) or sumr_75(5) or sumr_75(6) or sumr_75(7));
E(179)<=not ( sumr_76(0) or sumr_76(1) or sumr_76(2) or sumr_76(3) or sumr_76(4) or sumr_76(5) or sumr_76(6) or sumr_76(7));
E(178)<=not ( sumr_77(0) or sumr_77(1) or sumr_77(2) or sumr_77(3) or sumr_77(4) or sumr_77(5) or sumr_77(6) or sumr_77(7));
E(177)<=not ( sumr_78(0) or sumr_78(1) or sumr_78(2) or sumr_78(3) or sumr_78(4) or sumr_78(5) or sumr_78(6) or sumr_78(7));
E(176)<=not ( sumr_79(0) or sumr_79(1) or sumr_79(2) or sumr_79(3) or sumr_79(4) or sumr_79(5) or sumr_79(6) or sumr_79(7));
E(175)<=not ( sumr_80(0) or sumr_80(1) or sumr_80(2) or sumr_80(3) or sumr_80(4) or sumr_80(5) or sumr_80(6) or sumr_80(7));
E(174)<=not ( sumr_81(0) or sumr_81(1) or sumr_81(2) or sumr_81(3) or sumr_81(4) or sumr_81(5) or sumr_81(6) or sumr_81(7));
E(173)<=not ( sumr_82(0) or sumr_82(1) or sumr_82(2) or sumr_82(3) or sumr_82(4) or sumr_82(5) or sumr_82(6) or sumr_82(7));
E(172)<=not ( sumr_83(0) or sumr_83(1) or sumr_83(2) or sumr_83(3) or sumr_83(4) or sumr_83(5) or sumr_83(6) or sumr_83(7));
E(171)<=not ( sumr_84(0) or sumr_84(1) or sumr_84(2) or sumr_84(3) or sumr_84(4) or sumr_84(5) or sumr_84(6) or sumr_84(7));
E(170)<=not ( sumr_85(0) or sumr_85(1) or sumr_85(2) or sumr_85(3) or sumr_85(4) or sumr_85(5) or sumr_85(6) or sumr_85(7));
E(169)<=not ( sumr_86(0) or sumr_86(1) or sumr_86(2) or sumr_86(3) or sumr_86(4) or sumr_86(5) or sumr_86(6) or sumr_86(7));
E(168)<=not ( sumr_87(0) or sumr_87(1) or sumr_87(2) or sumr_87(3) or sumr_87(4) or sumr_87(5) or sumr_87(6) or sumr_87(7));
E(167)<=not ( sumr_88(0) or sumr_88(1) or sumr_88(2) or sumr_88(3) or sumr_88(4) or sumr_88(5) or sumr_88(6) or sumr_88(7));
E(166)<=not ( sumr_89(0) or sumr_89(1) or sumr_89(2) or sumr_89(3) or sumr_89(4) or sumr_89(5) or sumr_89(6) or sumr_89(7));
E(165)<=not ( sumr_90(0) or sumr_90(1) or sumr_90(2) or sumr_90(3) or sumr_90(4) or sumr_90(5) or sumr_90(6) or sumr_90(7));
E(164)<=not ( sumr_91(0) or sumr_91(1) or sumr_91(2) or sumr_91(3) or sumr_91(4) or sumr_91(5) or sumr_91(6) or sumr_91(7));
E(163)<=not ( sumr_92(0) or sumr_92(1) or sumr_92(2) or sumr_92(3) or sumr_92(4) or sumr_92(5) or sumr_92(6) or sumr_92(7));
E(162)<=not ( sumr_93(0) or sumr_93(1) or sumr_93(2) or sumr_93(3) or sumr_93(4) or sumr_93(5) or sumr_93(6) or sumr_93(7));
E(161)<=not ( sumr_94(0) or sumr_94(1) or sumr_94(2) or sumr_94(3) or sumr_94(4) or sumr_94(5) or sumr_94(6) or sumr_94(7));
E(160)<=not ( sumr_95(0) or sumr_95(1) or sumr_95(2) or sumr_95(3) or sumr_95(4) or sumr_95(5) or sumr_95(6) or sumr_95(7));
E(159)<=not ( sumr_96(0) or sumr_96(1) or sumr_96(2) or sumr_96(3) or sumr_96(4) or sumr_96(5) or sumr_96(6) or sumr_96(7));
E(158)<=not ( sumr_97(0) or sumr_97(1) or sumr_97(2) or sumr_97(3) or sumr_97(4) or sumr_97(5) or sumr_97(6) or sumr_97(7));
E(157)<=not ( sumr_98(0) or sumr_98(1) or sumr_98(2) or sumr_98(3) or sumr_98(4) or sumr_98(5) or sumr_98(6) or sumr_98(7));
E(156)<=not ( sumr_99(0) or sumr_99(1) or sumr_99(2) or sumr_99(3) or sumr_99(4) or sumr_99(5) or sumr_99(6) or sumr_99(7));
E(155)<=not ( sumr_100(0) or sumr_100(1) or sumr_100(2) or sumr_100(3) or sumr_100(4) or sumr_100(5) or sumr_100(6) or sumr_100(7));
E(154)<=not ( sumr_101(0) or sumr_101(1) or sumr_101(2) or sumr_101(3) or sumr_101(4) or sumr_101(5) or sumr_101(6) or sumr_101(7));
E(153)<=not ( sumr_102(0) or sumr_102(1) or sumr_102(2) or sumr_102(3) or sumr_102(4) or sumr_102(5) or sumr_102(6) or sumr_102(7));
E(152)<=not ( sumr_103(0) or sumr_103(1) or sumr_103(2) or sumr_103(3) or sumr_103(4) or sumr_103(5) or sumr_103(6) or sumr_103(7));
E(151)<=not ( sumr_104(0) or sumr_104(1) or sumr_104(2) or sumr_104(3) or sumr_104(4) or sumr_104(5) or sumr_104(6) or sumr_104(7));
E(150)<=not ( sumr_105(0) or sumr_105(1) or sumr_105(2) or sumr_105(3) or sumr_105(4) or sumr_105(5) or sumr_105(6) or sumr_105(7));
E(149)<=not ( sumr_106(0) or sumr_106(1) or sumr_106(2) or sumr_106(3) or sumr_106(4) or sumr_106(5) or sumr_106(6) or sumr_106(7));
E(148)<=not ( sumr_107(0) or sumr_107(1) or sumr_107(2) or sumr_107(3) or sumr_107(4) or sumr_107(5) or sumr_107(6) or sumr_107(7));
E(147)<=not ( sumr_108(0) or sumr_108(1) or sumr_108(2) or sumr_108(3) or sumr_108(4) or sumr_108(5) or sumr_108(6) or sumr_108(7));
E(146)<=not ( sumr_109(0) or sumr_109(1) or sumr_109(2) or sumr_109(3) or sumr_109(4) or sumr_109(5) or sumr_109(6) or sumr_109(7));
E(145)<=not ( sumr_110(0) or sumr_110(1) or sumr_110(2) or sumr_110(3) or sumr_110(4) or sumr_110(5) or sumr_110(6) or sumr_110(7));
E(144)<=not ( sumr_111(0) or sumr_111(1) or sumr_111(2) or sumr_111(3) or sumr_111(4) or sumr_111(5) or sumr_111(6) or sumr_111(7));
E(143)<=not ( sumr_112(0) or sumr_112(1) or sumr_112(2) or sumr_112(3) or sumr_112(4) or sumr_112(5) or sumr_112(6) or sumr_112(7));
E(142)<=not ( sumr_113(0) or sumr_113(1) or sumr_113(2) or sumr_113(3) or sumr_113(4) or sumr_113(5) or sumr_113(6) or sumr_113(7));
E(141)<=not ( sumr_114(0) or sumr_114(1) or sumr_114(2) or sumr_114(3) or sumr_114(4) or sumr_114(5) or sumr_114(6) or sumr_114(7));
E(140)<=not ( sumr_115(0) or sumr_115(1) or sumr_115(2) or sumr_115(3) or sumr_115(4) or sumr_115(5) or sumr_115(6) or sumr_115(7));
E(139)<=not ( sumr_116(0) or sumr_116(1) or sumr_116(2) or sumr_116(3) or sumr_116(4) or sumr_116(5) or sumr_116(6) or sumr_116(7));
E(138)<=not ( sumr_117(0) or sumr_117(1) or sumr_117(2) or sumr_117(3) or sumr_117(4) or sumr_117(5) or sumr_117(6) or sumr_117(7));
E(137)<=not ( sumr_118(0) or sumr_118(1) or sumr_118(2) or sumr_118(3) or sumr_118(4) or sumr_118(5) or sumr_118(6) or sumr_118(7));
E(136)<=not ( sumr_119(0) or sumr_119(1) or sumr_119(2) or sumr_119(3) or sumr_119(4) or sumr_119(5) or sumr_119(6) or sumr_119(7));
E(135)<=not ( sumr_120(0) or sumr_120(1) or sumr_120(2) or sumr_120(3) or sumr_120(4) or sumr_120(5) or sumr_120(6) or sumr_120(7));
E(134)<=not ( sumr_121(0) or sumr_121(1) or sumr_121(2) or sumr_121(3) or sumr_121(4) or sumr_121(5) or sumr_121(6) or sumr_121(7));
E(133)<=not ( sumr_122(0) or sumr_122(1) or sumr_122(2) or sumr_122(3) or sumr_122(4) or sumr_122(5) or sumr_122(6) or sumr_122(7));
E(132)<=not ( sumr_123(0) or sumr_123(1) or sumr_123(2) or sumr_123(3) or sumr_123(4) or sumr_123(5) or sumr_123(6) or sumr_123(7));
E(131)<=not ( sumr_124(0) or sumr_124(1) or sumr_124(2) or sumr_124(3) or sumr_124(4) or sumr_124(5) or sumr_124(6) or sumr_124(7));
E(130)<=not ( sumr_125(0) or sumr_125(1) or sumr_125(2) or sumr_125(3) or sumr_125(4) or sumr_125(5) or sumr_125(6) or sumr_125(7));
E(129)<=not ( sumr_126(0) or sumr_126(1) or sumr_126(2) or sumr_126(3) or sumr_126(4) or sumr_126(5) or sumr_126(6) or sumr_126(7));
E(128)<=not ( sumr_127(0) or sumr_127(1) or sumr_127(2) or sumr_127(3) or sumr_127(4) or sumr_127(5) or sumr_127(6) or sumr_127(7));
E(127)<=not ( sumr_128(0) or sumr_128(1) or sumr_128(2) or sumr_128(3) or sumr_128(4) or sumr_128(5) or sumr_128(6) or sumr_128(7));
E(126)<=not ( sumr_129(0) or sumr_129(1) or sumr_129(2) or sumr_129(3) or sumr_129(4) or sumr_129(5) or sumr_129(6) or sumr_129(7));
E(125)<=not ( sumr_130(0) or sumr_130(1) or sumr_130(2) or sumr_130(3) or sumr_130(4) or sumr_130(5) or sumr_130(6) or sumr_130(7));
E(124)<=not ( sumr_131(0) or sumr_131(1) or sumr_131(2) or sumr_131(3) or sumr_131(4) or sumr_131(5) or sumr_131(6) or sumr_131(7));
E(123)<=not ( sumr_132(0) or sumr_132(1) or sumr_132(2) or sumr_132(3) or sumr_132(4) or sumr_132(5) or sumr_132(6) or sumr_132(7));
E(122)<=not ( sumr_133(0) or sumr_133(1) or sumr_133(2) or sumr_133(3) or sumr_133(4) or sumr_133(5) or sumr_133(6) or sumr_133(7));
E(121)<=not ( sumr_134(0) or sumr_134(1) or sumr_134(2) or sumr_134(3) or sumr_134(4) or sumr_134(5) or sumr_134(6) or sumr_134(7));
E(120)<=not ( sumr_135(0) or sumr_135(1) or sumr_135(2) or sumr_135(3) or sumr_135(4) or sumr_135(5) or sumr_135(6) or sumr_135(7));
E(119)<=not ( sumr_136(0) or sumr_136(1) or sumr_136(2) or sumr_136(3) or sumr_136(4) or sumr_136(5) or sumr_136(6) or sumr_136(7));
E(118)<=not ( sumr_137(0) or sumr_137(1) or sumr_137(2) or sumr_137(3) or sumr_137(4) or sumr_137(5) or sumr_137(6) or sumr_137(7));
E(117)<=not ( sumr_138(0) or sumr_138(1) or sumr_138(2) or sumr_138(3) or sumr_138(4) or sumr_138(5) or sumr_138(6) or sumr_138(7));
E(116)<=not ( sumr_139(0) or sumr_139(1) or sumr_139(2) or sumr_139(3) or sumr_139(4) or sumr_139(5) or sumr_139(6) or sumr_139(7));
E(115)<=not ( sumr_140(0) or sumr_140(1) or sumr_140(2) or sumr_140(3) or sumr_140(4) or sumr_140(5) or sumr_140(6) or sumr_140(7));
E(114)<=not ( sumr_141(0) or sumr_141(1) or sumr_141(2) or sumr_141(3) or sumr_141(4) or sumr_141(5) or sumr_141(6) or sumr_141(7));
E(113)<=not ( sumr_142(0) or sumr_142(1) or sumr_142(2) or sumr_142(3) or sumr_142(4) or sumr_142(5) or sumr_142(6) or sumr_142(7));
E(112)<=not ( sumr_143(0) or sumr_143(1) or sumr_143(2) or sumr_143(3) or sumr_143(4) or sumr_143(5) or sumr_143(6) or sumr_143(7));
E(111)<=not ( sumr_144(0) or sumr_144(1) or sumr_144(2) or sumr_144(3) or sumr_144(4) or sumr_144(5) or sumr_144(6) or sumr_144(7));
E(110)<=not ( sumr_145(0) or sumr_145(1) or sumr_145(2) or sumr_145(3) or sumr_145(4) or sumr_145(5) or sumr_145(6) or sumr_145(7));
E(109)<=not ( sumr_146(0) or sumr_146(1) or sumr_146(2) or sumr_146(3) or sumr_146(4) or sumr_146(5) or sumr_146(6) or sumr_146(7));
E(108)<=not ( sumr_147(0) or sumr_147(1) or sumr_147(2) or sumr_147(3) or sumr_147(4) or sumr_147(5) or sumr_147(6) or sumr_147(7));
E(107)<=not ( sumr_148(0) or sumr_148(1) or sumr_148(2) or sumr_148(3) or sumr_148(4) or sumr_148(5) or sumr_148(6) or sumr_148(7));
E(106)<=not ( sumr_149(0) or sumr_149(1) or sumr_149(2) or sumr_149(3) or sumr_149(4) or sumr_149(5) or sumr_149(6) or sumr_149(7));
E(105)<=not ( sumr_150(0) or sumr_150(1) or sumr_150(2) or sumr_150(3) or sumr_150(4) or sumr_150(5) or sumr_150(6) or sumr_150(7));
E(104)<=not ( sumr_151(0) or sumr_151(1) or sumr_151(2) or sumr_151(3) or sumr_151(4) or sumr_151(5) or sumr_151(6) or sumr_151(7));
E(103)<=not ( sumr_152(0) or sumr_152(1) or sumr_152(2) or sumr_152(3) or sumr_152(4) or sumr_152(5) or sumr_152(6) or sumr_152(7));
E(102)<=not ( sumr_153(0) or sumr_153(1) or sumr_153(2) or sumr_153(3) or sumr_153(4) or sumr_153(5) or sumr_153(6) or sumr_153(7));
E(101)<=not ( sumr_154(0) or sumr_154(1) or sumr_154(2) or sumr_154(3) or sumr_154(4) or sumr_154(5) or sumr_154(6) or sumr_154(7));
E(100)<=not ( sumr_155(0) or sumr_155(1) or sumr_155(2) or sumr_155(3) or sumr_155(4) or sumr_155(5) or sumr_155(6) or sumr_155(7));
E(99)<=not ( sumr_156(0) or sumr_156(1) or sumr_156(2) or sumr_156(3) or sumr_156(4) or sumr_156(5) or sumr_156(6) or sumr_156(7));
E(98)<=not ( sumr_157(0) or sumr_157(1) or sumr_157(2) or sumr_157(3) or sumr_157(4) or sumr_157(5) or sumr_157(6) or sumr_157(7));
E(97)<=not ( sumr_158(0) or sumr_158(1) or sumr_158(2) or sumr_158(3) or sumr_158(4) or sumr_158(5) or sumr_158(6) or sumr_158(7));
E(96)<=not ( sumr_159(0) or sumr_159(1) or sumr_159(2) or sumr_159(3) or sumr_159(4) or sumr_159(5) or sumr_159(6) or sumr_159(7));
E(95)<=not ( sumr_160(0) or sumr_160(1) or sumr_160(2) or sumr_160(3) or sumr_160(4) or sumr_160(5) or sumr_160(6) or sumr_160(7));
E(94)<=not ( sumr_161(0) or sumr_161(1) or sumr_161(2) or sumr_161(3) or sumr_161(4) or sumr_161(5) or sumr_161(6) or sumr_161(7));
E(93)<=not ( sumr_162(0) or sumr_162(1) or sumr_162(2) or sumr_162(3) or sumr_162(4) or sumr_162(5) or sumr_162(6) or sumr_162(7));
E(92)<=not ( sumr_163(0) or sumr_163(1) or sumr_163(2) or sumr_163(3) or sumr_163(4) or sumr_163(5) or sumr_163(6) or sumr_163(7));
E(91)<=not ( sumr_164(0) or sumr_164(1) or sumr_164(2) or sumr_164(3) or sumr_164(4) or sumr_164(5) or sumr_164(6) or sumr_164(7));
E(90)<=not ( sumr_165(0) or sumr_165(1) or sumr_165(2) or sumr_165(3) or sumr_165(4) or sumr_165(5) or sumr_165(6) or sumr_165(7));
E(89)<=not ( sumr_166(0) or sumr_166(1) or sumr_166(2) or sumr_166(3) or sumr_166(4) or sumr_166(5) or sumr_166(6) or sumr_166(7));
E(88)<=not ( sumr_167(0) or sumr_167(1) or sumr_167(2) or sumr_167(3) or sumr_167(4) or sumr_167(5) or sumr_167(6) or sumr_167(7));
E(87)<=not ( sumr_168(0) or sumr_168(1) or sumr_168(2) or sumr_168(3) or sumr_168(4) or sumr_168(5) or sumr_168(6) or sumr_168(7));
E(86)<=not ( sumr_169(0) or sumr_169(1) or sumr_169(2) or sumr_169(3) or sumr_169(4) or sumr_169(5) or sumr_169(6) or sumr_169(7));
E(85)<=not ( sumr_170(0) or sumr_170(1) or sumr_170(2) or sumr_170(3) or sumr_170(4) or sumr_170(5) or sumr_170(6) or sumr_170(7));
E(84)<=not ( sumr_171(0) or sumr_171(1) or sumr_171(2) or sumr_171(3) or sumr_171(4) or sumr_171(5) or sumr_171(6) or sumr_171(7));
E(83)<=not ( sumr_172(0) or sumr_172(1) or sumr_172(2) or sumr_172(3) or sumr_172(4) or sumr_172(5) or sumr_172(6) or sumr_172(7));
E(82)<=not ( sumr_173(0) or sumr_173(1) or sumr_173(2) or sumr_173(3) or sumr_173(4) or sumr_173(5) or sumr_173(6) or sumr_173(7));
E(81)<=not ( sumr_174(0) or sumr_174(1) or sumr_174(2) or sumr_174(3) or sumr_174(4) or sumr_174(5) or sumr_174(6) or sumr_174(7));
E(80)<=not ( sumr_175(0) or sumr_175(1) or sumr_175(2) or sumr_175(3) or sumr_175(4) or sumr_175(5) or sumr_175(6) or sumr_175(7));
E(79)<=not ( sumr_176(0) or sumr_176(1) or sumr_176(2) or sumr_176(3) or sumr_176(4) or sumr_176(5) or sumr_176(6) or sumr_176(7));
E(78)<=not ( sumr_177(0) or sumr_177(1) or sumr_177(2) or sumr_177(3) or sumr_177(4) or sumr_177(5) or sumr_177(6) or sumr_177(7));
E(77)<=not ( sumr_178(0) or sumr_178(1) or sumr_178(2) or sumr_178(3) or sumr_178(4) or sumr_178(5) or sumr_178(6) or sumr_178(7));
E(76)<=not ( sumr_179(0) or sumr_179(1) or sumr_179(2) or sumr_179(3) or sumr_179(4) or sumr_179(5) or sumr_179(6) or sumr_179(7));
E(75)<=not ( sumr_180(0) or sumr_180(1) or sumr_180(2) or sumr_180(3) or sumr_180(4) or sumr_180(5) or sumr_180(6) or sumr_180(7));
E(74)<=not ( sumr_181(0) or sumr_181(1) or sumr_181(2) or sumr_181(3) or sumr_181(4) or sumr_181(5) or sumr_181(6) or sumr_181(7));
E(73)<=not ( sumr_182(0) or sumr_182(1) or sumr_182(2) or sumr_182(3) or sumr_182(4) or sumr_182(5) or sumr_182(6) or sumr_182(7));
E(72)<=not ( sumr_183(0) or sumr_183(1) or sumr_183(2) or sumr_183(3) or sumr_183(4) or sumr_183(5) or sumr_183(6) or sumr_183(7));
E(71)<=not ( sumr_184(0) or sumr_184(1) or sumr_184(2) or sumr_184(3) or sumr_184(4) or sumr_184(5) or sumr_184(6) or sumr_184(7));
E(70)<=not ( sumr_185(0) or sumr_185(1) or sumr_185(2) or sumr_185(3) or sumr_185(4) or sumr_185(5) or sumr_185(6) or sumr_185(7));
E(69)<=not ( sumr_186(0) or sumr_186(1) or sumr_186(2) or sumr_186(3) or sumr_186(4) or sumr_186(5) or sumr_186(6) or sumr_186(7));
E(68)<=not ( sumr_187(0) or sumr_187(1) or sumr_187(2) or sumr_187(3) or sumr_187(4) or sumr_187(5) or sumr_187(6) or sumr_187(7));
E(67)<=not ( sumr_188(0) or sumr_188(1) or sumr_188(2) or sumr_188(3) or sumr_188(4) or sumr_188(5) or sumr_188(6) or sumr_188(7));
E(66)<=not ( sumr_189(0) or sumr_189(1) or sumr_189(2) or sumr_189(3) or sumr_189(4) or sumr_189(5) or sumr_189(6) or sumr_189(7));
E(65)<=not ( sumr_190(0) or sumr_190(1) or sumr_190(2) or sumr_190(3) or sumr_190(4) or sumr_190(5) or sumr_190(6) or sumr_190(7));
E(64)<=not ( sumr_191(0) or sumr_191(1) or sumr_191(2) or sumr_191(3) or sumr_191(4) or sumr_191(5) or sumr_191(6) or sumr_191(7));
E(63)<=not ( sumr_192(0) or sumr_192(1) or sumr_192(2) or sumr_192(3) or sumr_192(4) or sumr_192(5) or sumr_192(6) or sumr_192(7));
E(62)<=not ( sumr_193(0) or sumr_193(1) or sumr_193(2) or sumr_193(3) or sumr_193(4) or sumr_193(5) or sumr_193(6) or sumr_193(7));
E(61)<=not ( sumr_194(0) or sumr_194(1) or sumr_194(2) or sumr_194(3) or sumr_194(4) or sumr_194(5) or sumr_194(6) or sumr_194(7));
E(60)<=not ( sumr_195(0) or sumr_195(1) or sumr_195(2) or sumr_195(3) or sumr_195(4) or sumr_195(5) or sumr_195(6) or sumr_195(7));
E(59)<=not ( sumr_196(0) or sumr_196(1) or sumr_196(2) or sumr_196(3) or sumr_196(4) or sumr_196(5) or sumr_196(6) or sumr_196(7));
E(58)<=not ( sumr_197(0) or sumr_197(1) or sumr_197(2) or sumr_197(3) or sumr_197(4) or sumr_197(5) or sumr_197(6) or sumr_197(7));
E(57)<=not ( sumr_198(0) or sumr_198(1) or sumr_198(2) or sumr_198(3) or sumr_198(4) or sumr_198(5) or sumr_198(6) or sumr_198(7));
E(56)<=not ( sumr_199(0) or sumr_199(1) or sumr_199(2) or sumr_199(3) or sumr_199(4) or sumr_199(5) or sumr_199(6) or sumr_199(7));
E(55)<=not ( sumr_200(0) or sumr_200(1) or sumr_200(2) or sumr_200(3) or sumr_200(4) or sumr_200(5) or sumr_200(6) or sumr_200(7));
E(54)<=not ( sumr_201(0) or sumr_201(1) or sumr_201(2) or sumr_201(3) or sumr_201(4) or sumr_201(5) or sumr_201(6) or sumr_201(7));
E(53)<=not ( sumr_202(0) or sumr_202(1) or sumr_202(2) or sumr_202(3) or sumr_202(4) or sumr_202(5) or sumr_202(6) or sumr_202(7));
E(52)<=not ( sumr_203(0) or sumr_203(1) or sumr_203(2) or sumr_203(3) or sumr_203(4) or sumr_203(5) or sumr_203(6) or sumr_203(7));
E(51)<=not ( sumr_204(0) or sumr_204(1) or sumr_204(2) or sumr_204(3) or sumr_204(4) or sumr_204(5) or sumr_204(6) or sumr_204(7));
E(50)<=not ( sumr_205(0) or sumr_205(1) or sumr_205(2) or sumr_205(3) or sumr_205(4) or sumr_205(5) or sumr_205(6) or sumr_205(7));
E(49)<=not ( sumr_206(0) or sumr_206(1) or sumr_206(2) or sumr_206(3) or sumr_206(4) or sumr_206(5) or sumr_206(6) or sumr_206(7));
E(48)<=not ( sumr_207(0) or sumr_207(1) or sumr_207(2) or sumr_207(3) or sumr_207(4) or sumr_207(5) or sumr_207(6) or sumr_207(7));
E(47)<=not ( sumr_208(0) or sumr_208(1) or sumr_208(2) or sumr_208(3) or sumr_208(4) or sumr_208(5) or sumr_208(6) or sumr_208(7));
E(46)<=not ( sumr_209(0) or sumr_209(1) or sumr_209(2) or sumr_209(3) or sumr_209(4) or sumr_209(5) or sumr_209(6) or sumr_209(7));
E(45)<=not ( sumr_210(0) or sumr_210(1) or sumr_210(2) or sumr_210(3) or sumr_210(4) or sumr_210(5) or sumr_210(6) or sumr_210(7));
E(44)<=not ( sumr_211(0) or sumr_211(1) or sumr_211(2) or sumr_211(3) or sumr_211(4) or sumr_211(5) or sumr_211(6) or sumr_211(7));
E(43)<=not ( sumr_212(0) or sumr_212(1) or sumr_212(2) or sumr_212(3) or sumr_212(4) or sumr_212(5) or sumr_212(6) or sumr_212(7));
E(42)<=not ( sumr_213(0) or sumr_213(1) or sumr_213(2) or sumr_213(3) or sumr_213(4) or sumr_213(5) or sumr_213(6) or sumr_213(7));
E(41)<=not ( sumr_214(0) or sumr_214(1) or sumr_214(2) or sumr_214(3) or sumr_214(4) or sumr_214(5) or sumr_214(6) or sumr_214(7));
E(40)<=not ( sumr_215(0) or sumr_215(1) or sumr_215(2) or sumr_215(3) or sumr_215(4) or sumr_215(5) or sumr_215(6) or sumr_215(7));
E(39)<=not ( sumr_216(0) or sumr_216(1) or sumr_216(2) or sumr_216(3) or sumr_216(4) or sumr_216(5) or sumr_216(6) or sumr_216(7));
E(38)<=not ( sumr_217(0) or sumr_217(1) or sumr_217(2) or sumr_217(3) or sumr_217(4) or sumr_217(5) or sumr_217(6) or sumr_217(7));
E(37)<=not ( sumr_218(0) or sumr_218(1) or sumr_218(2) or sumr_218(3) or sumr_218(4) or sumr_218(5) or sumr_218(6) or sumr_218(7));
E(36)<=not ( sumr_219(0) or sumr_219(1) or sumr_219(2) or sumr_219(3) or sumr_219(4) or sumr_219(5) or sumr_219(6) or sumr_219(7));
E(35)<=not ( sumr_220(0) or sumr_220(1) or sumr_220(2) or sumr_220(3) or sumr_220(4) or sumr_220(5) or sumr_220(6) or sumr_220(7));
E(34)<=not ( sumr_221(0) or sumr_221(1) or sumr_221(2) or sumr_221(3) or sumr_221(4) or sumr_221(5) or sumr_221(6) or sumr_221(7));
E(33)<=not ( sumr_222(0) or sumr_222(1) or sumr_222(2) or sumr_222(3) or sumr_222(4) or sumr_222(5) or sumr_222(6) or sumr_222(7));
E(32)<=not ( sumr_223(0) or sumr_223(1) or sumr_223(2) or sumr_223(3) or sumr_223(4) or sumr_223(5) or sumr_223(6) or sumr_223(7));
E(31)<=not ( sumr_224(0) or sumr_224(1) or sumr_224(2) or sumr_224(3) or sumr_224(4) or sumr_224(5) or sumr_224(6) or sumr_224(7));
E(30)<=not ( sumr_225(0) or sumr_225(1) or sumr_225(2) or sumr_225(3) or sumr_225(4) or sumr_225(5) or sumr_225(6) or sumr_225(7));
E(29)<=not ( sumr_226(0) or sumr_226(1) or sumr_226(2) or sumr_226(3) or sumr_226(4) or sumr_226(5) or sumr_226(6) or sumr_226(7));
E(28)<=not ( sumr_227(0) or sumr_227(1) or sumr_227(2) or sumr_227(3) or sumr_227(4) or sumr_227(5) or sumr_227(6) or sumr_227(7));
E(27)<=not ( sumr_228(0) or sumr_228(1) or sumr_228(2) or sumr_228(3) or sumr_228(4) or sumr_228(5) or sumr_228(6) or sumr_228(7));
E(26)<=not ( sumr_229(0) or sumr_229(1) or sumr_229(2) or sumr_229(3) or sumr_229(4) or sumr_229(5) or sumr_229(6) or sumr_229(7));
E(25)<=not ( sumr_230(0) or sumr_230(1) or sumr_230(2) or sumr_230(3) or sumr_230(4) or sumr_230(5) or sumr_230(6) or sumr_230(7));
E(24)<=not ( sumr_231(0) or sumr_231(1) or sumr_231(2) or sumr_231(3) or sumr_231(4) or sumr_231(5) or sumr_231(6) or sumr_231(7));
E(23)<=not ( sumr_232(0) or sumr_232(1) or sumr_232(2) or sumr_232(3) or sumr_232(4) or sumr_232(5) or sumr_232(6) or sumr_232(7));
E(22)<=not ( sumr_233(0) or sumr_233(1) or sumr_233(2) or sumr_233(3) or sumr_233(4) or sumr_233(5) or sumr_233(6) or sumr_233(7));
E(21)<=not ( sumr_234(0) or sumr_234(1) or sumr_234(2) or sumr_234(3) or sumr_234(4) or sumr_234(5) or sumr_234(6) or sumr_234(7));
E(20)<=not ( sumr_235(0) or sumr_235(1) or sumr_235(2) or sumr_235(3) or sumr_235(4) or sumr_235(5) or sumr_235(6) or sumr_235(7));
E(19)<=not ( sumr_236(0) or sumr_236(1) or sumr_236(2) or sumr_236(3) or sumr_236(4) or sumr_236(5) or sumr_236(6) or sumr_236(7));
E(18)<=not ( sumr_237(0) or sumr_237(1) or sumr_237(2) or sumr_237(3) or sumr_237(4) or sumr_237(5) or sumr_237(6) or sumr_237(7));
E(17)<=not ( sumr_238(0) or sumr_238(1) or sumr_238(2) or sumr_238(3) or sumr_238(4) or sumr_238(5) or sumr_238(6) or sumr_238(7));
E(16)<=not ( sumr_239(0) or sumr_239(1) or sumr_239(2) or sumr_239(3) or sumr_239(4) or sumr_239(5) or sumr_239(6) or sumr_239(7));
E(15)<=not ( sumr_240(0) or sumr_240(1) or sumr_240(2) or sumr_240(3) or sumr_240(4) or sumr_240(5) or sumr_240(6) or sumr_240(7));
E(14)<=not ( sumr_241(0) or sumr_241(1) or sumr_241(2) or sumr_241(3) or sumr_241(4) or sumr_241(5) or sumr_241(6) or sumr_241(7));
E(13)<=not ( sumr_242(0) or sumr_242(1) or sumr_242(2) or sumr_242(3) or sumr_242(4) or sumr_242(5) or sumr_242(6) or sumr_242(7));
E(12)<=not ( sumr_243(0) or sumr_243(1) or sumr_243(2) or sumr_243(3) or sumr_243(4) or sumr_243(5) or sumr_243(6) or sumr_243(7));
E(11)<=not ( sumr_244(0) or sumr_244(1) or sumr_244(2) or sumr_244(3) or sumr_244(4) or sumr_244(5) or sumr_244(6) or sumr_244(7));
E(10)<=not ( sumr_245(0) or sumr_245(1) or sumr_245(2) or sumr_245(3) or sumr_245(4) or sumr_245(5) or sumr_245(6) or sumr_245(7));
E(9)<=not ( sumr_246(0) or sumr_246(1) or sumr_246(2) or sumr_246(3) or sumr_246(4) or sumr_246(5) or sumr_246(6) or sumr_246(7));
E(8)<=not ( sumr_247(0) or sumr_247(1) or sumr_247(2) or sumr_247(3) or sumr_247(4) or sumr_247(5) or sumr_247(6) or sumr_247(7));
E(7)<=not ( sumr_248(0) or sumr_248(1) or sumr_248(2) or sumr_248(3) or sumr_248(4) or sumr_248(5) or sumr_248(6) or sumr_248(7));
E(6)<=not ( sumr_249(0) or sumr_249(1) or sumr_249(2) or sumr_249(3) or sumr_249(4) or sumr_249(5) or sumr_249(6) or sumr_249(7));
E(5)<=not ( sumr_250(0) or sumr_250(1) or sumr_250(2) or sumr_250(3) or sumr_250(4) or sumr_250(5) or sumr_250(6) or sumr_250(7));
E(4)<=not ( sumr_251(0) or sumr_251(1) or sumr_251(2) or sumr_251(3) or sumr_251(4) or sumr_251(5) or sumr_251(6) or sumr_251(7));
E(3)<=not ( sumr_252(0) or sumr_252(1) or sumr_252(2) or sumr_252(3) or sumr_252(4) or sumr_252(5) or sumr_252(6) or sumr_252(7));
E(2)<=not ( sumr_253(0) or sumr_253(1) or sumr_253(2) or sumr_253(3) or sumr_253(4) or sumr_253(5) or sumr_253(6) or sumr_253(7));
E(1)<=not ( sumr_254(0) or sumr_254(1) or sumr_254(2) or sumr_254(3) or sumr_254(4) or sumr_254(5) or sumr_254(6) or sumr_254(7));
E(0)<=not ( sumr_255(0) or sumr_255(1) or sumr_255(2) or sumr_255(3) or sumr_255(4) or sumr_255(5) or sumr_255(6) or sumr_255(7));
end arch;
