----------------------------------------------------------------------------------
    -- Company:  Chalmers
    -- Engineer: Fredrik Åkerlund
    -- 
    -- Create Date: Mon Jul 24 13:30:05 2017

    -- Design Name: 
    -- Module Name: word_expander_64IN_to_493OUT - arch_word_expander_64IN_to_493OUT
    -- Project Name: 
    -- Target Devices: 
    -- Tool Versions: 
    -- Description: 
    -- 
    -- Dependencies: 
    -- 
    -- Revision:
    -- Revision 0.01 - File Created
    -- Additional Comments:
    -- 
    ----------------------------------------------------------------------------------


    library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;

    -- Uncomment the following library declaration if using
    -- arithmetic functions with Signed or Unsigned values
    use IEEE.NUMERIC_STD.ALL;

    -- Uncomment the following library declaration if instantiating
    -- any Xilinx leaf cells in this code.
    --library UNISIM;
    --use UNISIM.VComponents.all;
    entity word_expander_64IN_to_493OUT is

    generic(
        IN_WIDTH  : integer := 64;
        OUT_WIDTH : integer := 493
    );
    port(
        user_clk  : in  std_logic;       
        reset_in  : in  std_logic;
        enable_in : in  std_logic;

        in_rdy    : in  std_logic;
        data_in   : in  std_logic_vector(IN_WIDTH-1 downto 0);

        buf_out   : out std_logic_vector(OUT_WIDTH-1 downto 0);
        out_rdy   : out std_logic

        );
    end word_expander_64IN_to_493OUT;
architecture arch_word_expander_64IN_to_493OUT of word_expander_64IN_to_493OUT is

        constant BUF_WIDTH : integer := (OUT_WIDTH + IN_WIDTH);

        signal buf_input_r  : std_logic_vector(BUF_WIDTH-1 downto 0);
        signal buf_output_r : std_logic_vector(OUT_WIDTH-1 downto 0);
        signal out_rdy_r    : std_logic;

        signal bits_in_buffer : integer range 0 to BUF_WIDTH;

    begin

    output_reg_process:
    process(reset_in, user_clk, enable_in)
    begin
        if reset_in = '0' then
            buf_out <= (others=>'0');
            out_rdy <= '0';
        elsif rising_edge(user_clk) then
            if enable_in = '1' then
                buf_out <= buf_output_r;
                out_rdy <= out_rdy_r;
            end if;
        end if;
    end process;


    the_buffing_process:
    process(reset_in, user_clk, in_rdy, enable_in)
    begin
        if reset_in = '0' then

            buf_input_r  <= (others=>'0');
            buf_output_r <= (others=>'0');

            bits_in_buffer <= 0;

            out_rdy_r <= '0';

        elsif rising_edge(user_clk) then
            if in_rdy = '1' and enable_in = '1' then
            if bits_in_buffer >= 429 then
                out_rdy_r <= '1';
                case bits_in_buffer is
                    when 429 =>
                        buf_output_r(428 downto 0)   <= buf_input_r(428 downto 0);
                        buf_output_r(492 downto 429) <= data_in(63 downto 0);
                        buf_input_r                  <= (others=>'0');
                        bits_in_buffer               <= 0;
                    when 430 =>
                        buf_output_r(429 downto 0)   <= buf_input_r(429 downto 0);
                        buf_output_r(492 downto 430) <= data_in(62 downto 0);
                        buf_input_r (0 downto 0)     <= data_in(63 downto 63);
                        bits_in_buffer               <= 1;
                    when 431 =>
                        buf_output_r(430 downto 0)   <= buf_input_r(430 downto 0);
                        buf_output_r(492 downto 431) <= data_in(61 downto 0);
                        buf_input_r (1 downto 0)     <= data_in(63 downto 62);
                        bits_in_buffer               <= 2;
                    when 432 =>
                        buf_output_r(431 downto 0)   <= buf_input_r(431 downto 0);
                        buf_output_r(492 downto 432) <= data_in(60 downto 0);
                        buf_input_r (2 downto 0)     <= data_in(63 downto 61);
                        bits_in_buffer               <= 3;
                    when 433 =>
                        buf_output_r(432 downto 0)   <= buf_input_r(432 downto 0);
                        buf_output_r(492 downto 433) <= data_in(59 downto 0);
                        buf_input_r (3 downto 0)     <= data_in(63 downto 60);
                        bits_in_buffer               <= 4;
                    when 434 =>
                        buf_output_r(433 downto 0)   <= buf_input_r(433 downto 0);
                        buf_output_r(492 downto 434) <= data_in(58 downto 0);
                        buf_input_r (4 downto 0)     <= data_in(63 downto 59);
                        bits_in_buffer               <= 5;
                    when 435 =>
                        buf_output_r(434 downto 0)   <= buf_input_r(434 downto 0);
                        buf_output_r(492 downto 435) <= data_in(57 downto 0);
                        buf_input_r (5 downto 0)     <= data_in(63 downto 58);
                        bits_in_buffer               <= 6;
                    when 436 =>
                        buf_output_r(435 downto 0)   <= buf_input_r(435 downto 0);
                        buf_output_r(492 downto 436) <= data_in(56 downto 0);
                        buf_input_r (6 downto 0)     <= data_in(63 downto 57);
                        bits_in_buffer               <= 7;
                    when 437 =>
                        buf_output_r(436 downto 0)   <= buf_input_r(436 downto 0);
                        buf_output_r(492 downto 437) <= data_in(55 downto 0);
                        buf_input_r (7 downto 0)     <= data_in(63 downto 56);
                        bits_in_buffer               <= 8;
                    when 438 =>
                        buf_output_r(437 downto 0)   <= buf_input_r(437 downto 0);
                        buf_output_r(492 downto 438) <= data_in(54 downto 0);
                        buf_input_r (8 downto 0)     <= data_in(63 downto 55);
                        bits_in_buffer               <= 9;
                    when 439 =>
                        buf_output_r(438 downto 0)   <= buf_input_r(438 downto 0);
                        buf_output_r(492 downto 439) <= data_in(53 downto 0);
                        buf_input_r (9 downto 0)     <= data_in(63 downto 54);
                        bits_in_buffer               <= 10;
                    when 440 =>
                        buf_output_r(439 downto 0)   <= buf_input_r(439 downto 0);
                        buf_output_r(492 downto 440) <= data_in(52 downto 0);
                        buf_input_r (10 downto 0)    <= data_in(63 downto 53);
                        bits_in_buffer               <= 11;
                    when 441 =>
                        buf_output_r(440 downto 0)   <= buf_input_r(440 downto 0);
                        buf_output_r(492 downto 441) <= data_in(51 downto 0);
                        buf_input_r (11 downto 0)    <= data_in(63 downto 52);
                        bits_in_buffer               <= 12;
                    when 442 =>
                        buf_output_r(441 downto 0)   <= buf_input_r(441 downto 0);
                        buf_output_r(492 downto 442) <= data_in(50 downto 0);
                        buf_input_r (12 downto 0)    <= data_in(63 downto 51);
                        bits_in_buffer               <= 13;
                    when 443 =>
                        buf_output_r(442 downto 0)   <= buf_input_r(442 downto 0);
                        buf_output_r(492 downto 443) <= data_in(49 downto 0);
                        buf_input_r (13 downto 0)    <= data_in(63 downto 50);
                        bits_in_buffer               <= 14;
                    when 444 =>
                        buf_output_r(443 downto 0)   <= buf_input_r(443 downto 0);
                        buf_output_r(492 downto 444) <= data_in(48 downto 0);
                        buf_input_r (14 downto 0)    <= data_in(63 downto 49);
                        bits_in_buffer               <= 15;
                    when 445 =>
                        buf_output_r(444 downto 0)   <= buf_input_r(444 downto 0);
                        buf_output_r(492 downto 445) <= data_in(47 downto 0);
                        buf_input_r (15 downto 0)    <= data_in(63 downto 48);
                        bits_in_buffer               <= 16;
                    when 446 =>
                        buf_output_r(445 downto 0)   <= buf_input_r(445 downto 0);
                        buf_output_r(492 downto 446) <= data_in(46 downto 0);
                        buf_input_r (16 downto 0)    <= data_in(63 downto 47);
                        bits_in_buffer               <= 17;
                    when 447 =>
                        buf_output_r(446 downto 0)   <= buf_input_r(446 downto 0);
                        buf_output_r(492 downto 447) <= data_in(45 downto 0);
                        buf_input_r (17 downto 0)    <= data_in(63 downto 46);
                        bits_in_buffer               <= 18;
                    when 448 =>
                        buf_output_r(447 downto 0)   <= buf_input_r(447 downto 0);
                        buf_output_r(492 downto 448) <= data_in(44 downto 0);
                        buf_input_r (18 downto 0)    <= data_in(63 downto 45);
                        bits_in_buffer               <= 19;
                    when 449 =>
                        buf_output_r(448 downto 0)   <= buf_input_r(448 downto 0);
                        buf_output_r(492 downto 449) <= data_in(43 downto 0);
                        buf_input_r (19 downto 0)    <= data_in(63 downto 44);
                        bits_in_buffer               <= 20;
                    when 450 =>
                        buf_output_r(449 downto 0)   <= buf_input_r(449 downto 0);
                        buf_output_r(492 downto 450) <= data_in(42 downto 0);
                        buf_input_r (20 downto 0)    <= data_in(63 downto 43);
                        bits_in_buffer               <= 21;
                    when 451 =>
                        buf_output_r(450 downto 0)   <= buf_input_r(450 downto 0);
                        buf_output_r(492 downto 451) <= data_in(41 downto 0);
                        buf_input_r (21 downto 0)    <= data_in(63 downto 42);
                        bits_in_buffer               <= 22;
                    when 452 =>
                        buf_output_r(451 downto 0)   <= buf_input_r(451 downto 0);
                        buf_output_r(492 downto 452) <= data_in(40 downto 0);
                        buf_input_r (22 downto 0)    <= data_in(63 downto 41);
                        bits_in_buffer               <= 23;
                    when 453 =>
                        buf_output_r(452 downto 0)   <= buf_input_r(452 downto 0);
                        buf_output_r(492 downto 453) <= data_in(39 downto 0);
                        buf_input_r (23 downto 0)    <= data_in(63 downto 40);
                        bits_in_buffer               <= 24;
                    when 454 =>
                        buf_output_r(453 downto 0)   <= buf_input_r(453 downto 0);
                        buf_output_r(492 downto 454) <= data_in(38 downto 0);
                        buf_input_r (24 downto 0)    <= data_in(63 downto 39);
                        bits_in_buffer               <= 25;
                    when 455 =>
                        buf_output_r(454 downto 0)   <= buf_input_r(454 downto 0);
                        buf_output_r(492 downto 455) <= data_in(37 downto 0);
                        buf_input_r (25 downto 0)    <= data_in(63 downto 38);
                        bits_in_buffer               <= 26;
                    when 456 =>
                        buf_output_r(455 downto 0)   <= buf_input_r(455 downto 0);
                        buf_output_r(492 downto 456) <= data_in(36 downto 0);
                        buf_input_r (26 downto 0)    <= data_in(63 downto 37);
                        bits_in_buffer               <= 27;
                    when 457 =>
                        buf_output_r(456 downto 0)   <= buf_input_r(456 downto 0);
                        buf_output_r(492 downto 457) <= data_in(35 downto 0);
                        buf_input_r (27 downto 0)    <= data_in(63 downto 36);
                        bits_in_buffer               <= 28;
                    when 458 =>
                        buf_output_r(457 downto 0)   <= buf_input_r(457 downto 0);
                        buf_output_r(492 downto 458) <= data_in(34 downto 0);
                        buf_input_r (28 downto 0)    <= data_in(63 downto 35);
                        bits_in_buffer               <= 29;
                    when 459 =>
                        buf_output_r(458 downto 0)   <= buf_input_r(458 downto 0);
                        buf_output_r(492 downto 459) <= data_in(33 downto 0);
                        buf_input_r (29 downto 0)    <= data_in(63 downto 34);
                        bits_in_buffer               <= 30;
                    when 460 =>
                        buf_output_r(459 downto 0)   <= buf_input_r(459 downto 0);
                        buf_output_r(492 downto 460) <= data_in(32 downto 0);
                        buf_input_r (30 downto 0)    <= data_in(63 downto 33);
                        bits_in_buffer               <= 31;
                    when 461 =>
                        buf_output_r(460 downto 0)   <= buf_input_r(460 downto 0);
                        buf_output_r(492 downto 461) <= data_in(31 downto 0);
                        buf_input_r (31 downto 0)    <= data_in(63 downto 32);
                        bits_in_buffer               <= 32;
                    when 462 =>
                        buf_output_r(461 downto 0)   <= buf_input_r(461 downto 0);
                        buf_output_r(492 downto 462) <= data_in(30 downto 0);
                        buf_input_r (32 downto 0)    <= data_in(63 downto 31);
                        bits_in_buffer               <= 33;
                    when 463 =>
                        buf_output_r(462 downto 0)   <= buf_input_r(462 downto 0);
                        buf_output_r(492 downto 463) <= data_in(29 downto 0);
                        buf_input_r (33 downto 0)    <= data_in(63 downto 30);
                        bits_in_buffer               <= 34;
                    when 464 =>
                        buf_output_r(463 downto 0)   <= buf_input_r(463 downto 0);
                        buf_output_r(492 downto 464) <= data_in(28 downto 0);
                        buf_input_r (34 downto 0)    <= data_in(63 downto 29);
                        bits_in_buffer               <= 35;
                    when 465 =>
                        buf_output_r(464 downto 0)   <= buf_input_r(464 downto 0);
                        buf_output_r(492 downto 465) <= data_in(27 downto 0);
                        buf_input_r (35 downto 0)    <= data_in(63 downto 28);
                        bits_in_buffer               <= 36;
                    when 466 =>
                        buf_output_r(465 downto 0)   <= buf_input_r(465 downto 0);
                        buf_output_r(492 downto 466) <= data_in(26 downto 0);
                        buf_input_r (36 downto 0)    <= data_in(63 downto 27);
                        bits_in_buffer               <= 37;
                    when 467 =>
                        buf_output_r(466 downto 0)   <= buf_input_r(466 downto 0);
                        buf_output_r(492 downto 467) <= data_in(25 downto 0);
                        buf_input_r (37 downto 0)    <= data_in(63 downto 26);
                        bits_in_buffer               <= 38;
                    when 468 =>
                        buf_output_r(467 downto 0)   <= buf_input_r(467 downto 0);
                        buf_output_r(492 downto 468) <= data_in(24 downto 0);
                        buf_input_r (38 downto 0)    <= data_in(63 downto 25);
                        bits_in_buffer               <= 39;
                    when 469 =>
                        buf_output_r(468 downto 0)   <= buf_input_r(468 downto 0);
                        buf_output_r(492 downto 469) <= data_in(23 downto 0);
                        buf_input_r (39 downto 0)    <= data_in(63 downto 24);
                        bits_in_buffer               <= 40;
                    when 470 =>
                        buf_output_r(469 downto 0)   <= buf_input_r(469 downto 0);
                        buf_output_r(492 downto 470) <= data_in(22 downto 0);
                        buf_input_r (40 downto 0)    <= data_in(63 downto 23);
                        bits_in_buffer               <= 41;
                    when 471 =>
                        buf_output_r(470 downto 0)   <= buf_input_r(470 downto 0);
                        buf_output_r(492 downto 471) <= data_in(21 downto 0);
                        buf_input_r (41 downto 0)    <= data_in(63 downto 22);
                        bits_in_buffer               <= 42;
                    when 472 =>
                        buf_output_r(471 downto 0)   <= buf_input_r(471 downto 0);
                        buf_output_r(492 downto 472) <= data_in(20 downto 0);
                        buf_input_r (42 downto 0)    <= data_in(63 downto 21);
                        bits_in_buffer               <= 43;
                    when 473 =>
                        buf_output_r(472 downto 0)   <= buf_input_r(472 downto 0);
                        buf_output_r(492 downto 473) <= data_in(19 downto 0);
                        buf_input_r (43 downto 0)    <= data_in(63 downto 20);
                        bits_in_buffer               <= 44;
                    when 474 =>
                        buf_output_r(473 downto 0)   <= buf_input_r(473 downto 0);
                        buf_output_r(492 downto 474) <= data_in(18 downto 0);
                        buf_input_r (44 downto 0)    <= data_in(63 downto 19);
                        bits_in_buffer               <= 45;
                    when 475 =>
                        buf_output_r(474 downto 0)   <= buf_input_r(474 downto 0);
                        buf_output_r(492 downto 475) <= data_in(17 downto 0);
                        buf_input_r (45 downto 0)    <= data_in(63 downto 18);
                        bits_in_buffer               <= 46;
                    when 476 =>
                        buf_output_r(475 downto 0)   <= buf_input_r(475 downto 0);
                        buf_output_r(492 downto 476) <= data_in(16 downto 0);
                        buf_input_r (46 downto 0)    <= data_in(63 downto 17);
                        bits_in_buffer               <= 47;
                    when 477 =>
                        buf_output_r(476 downto 0)   <= buf_input_r(476 downto 0);
                        buf_output_r(492 downto 477) <= data_in(15 downto 0);
                        buf_input_r (47 downto 0)    <= data_in(63 downto 16);
                        bits_in_buffer               <= 48;
                    when 478 =>
                        buf_output_r(477 downto 0)   <= buf_input_r(477 downto 0);
                        buf_output_r(492 downto 478) <= data_in(14 downto 0);
                        buf_input_r (48 downto 0)    <= data_in(63 downto 15);
                        bits_in_buffer               <= 49;
                    when 479 =>
                        buf_output_r(478 downto 0)   <= buf_input_r(478 downto 0);
                        buf_output_r(492 downto 479) <= data_in(13 downto 0);
                        buf_input_r (49 downto 0)    <= data_in(63 downto 14);
                        bits_in_buffer               <= 50;
                    when 480 =>
                        buf_output_r(479 downto 0)   <= buf_input_r(479 downto 0);
                        buf_output_r(492 downto 480) <= data_in(12 downto 0);
                        buf_input_r (50 downto 0)    <= data_in(63 downto 13);
                        bits_in_buffer               <= 51;
                    when 481 =>
                        buf_output_r(480 downto 0)   <= buf_input_r(480 downto 0);
                        buf_output_r(492 downto 481) <= data_in(11 downto 0);
                        buf_input_r (51 downto 0)    <= data_in(63 downto 12);
                        bits_in_buffer               <= 52;
                    when 482 =>
                        buf_output_r(481 downto 0)   <= buf_input_r(481 downto 0);
                        buf_output_r(492 downto 482) <= data_in(10 downto 0);
                        buf_input_r (52 downto 0)    <= data_in(63 downto 11);
                        bits_in_buffer               <= 53;
                    when 483 =>
                        buf_output_r(482 downto 0)   <= buf_input_r(482 downto 0);
                        buf_output_r(492 downto 483) <= data_in(9 downto 0);
                        buf_input_r (53 downto 0)    <= data_in(63 downto 10);
                        bits_in_buffer               <= 54;
                    when 484 =>
                        buf_output_r(483 downto 0)   <= buf_input_r(483 downto 0);
                        buf_output_r(492 downto 484) <= data_in(8 downto 0);
                        buf_input_r (54 downto 0)    <= data_in(63 downto 9);
                        bits_in_buffer               <= 55;
                    when 485 =>
                        buf_output_r(484 downto 0)   <= buf_input_r(484 downto 0);
                        buf_output_r(492 downto 485) <= data_in(7 downto 0);
                        buf_input_r (55 downto 0)    <= data_in(63 downto 8);
                        bits_in_buffer               <= 56;
                    when 486 =>
                        buf_output_r(485 downto 0)   <= buf_input_r(485 downto 0);
                        buf_output_r(492 downto 486) <= data_in(6 downto 0);
                        buf_input_r (56 downto 0)    <= data_in(63 downto 7);
                        bits_in_buffer               <= 57;
                    when 487 =>
                        buf_output_r(486 downto 0)   <= buf_input_r(486 downto 0);
                        buf_output_r(492 downto 487) <= data_in(5 downto 0);
                        buf_input_r (57 downto 0)    <= data_in(63 downto 6);
                        bits_in_buffer               <= 58;
                    when 488 =>
                        buf_output_r(487 downto 0)   <= buf_input_r(487 downto 0);
                        buf_output_r(492 downto 488) <= data_in(4 downto 0);
                        buf_input_r (58 downto 0)    <= data_in(63 downto 5);
                        bits_in_buffer               <= 59;
                    when 489 =>
                        buf_output_r(488 downto 0)   <= buf_input_r(488 downto 0);
                        buf_output_r(492 downto 489) <= data_in(3 downto 0);
                        buf_input_r (59 downto 0)    <= data_in(63 downto 4);
                        bits_in_buffer               <= 60;
                    when 490 =>
                        buf_output_r(489 downto 0)   <= buf_input_r(489 downto 0);
                        buf_output_r(492 downto 490) <= data_in(2 downto 0);
                        buf_input_r (60 downto 0)    <= data_in(63 downto 3);
                        bits_in_buffer               <= 61;
                    when 491 =>
                        buf_output_r(490 downto 0)   <= buf_input_r(490 downto 0);
                        buf_output_r(492 downto 491) <= data_in(1 downto 0);
                        buf_input_r (61 downto 0)    <= data_in(63 downto 2);
                        bits_in_buffer               <= 62;
                    when 492 =>
                        buf_output_r(491 downto 0)   <= buf_input_r(491 downto 0);
                        buf_output_r(492 downto 492) <= data_in(0 downto 0);
                        buf_input_r (62 downto 0)    <= data_in(63 downto 1);
                        bits_in_buffer               <= 63;
                    when others =>
                end case;
            else
                out_rdy_r <= '0';
                case bits_in_buffer is
                    when 0 =>
                        buf_input_r (63 downto 0)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 64;
                    when 1 =>
                        buf_input_r (64 downto 1)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 65;
                    when 2 =>
                        buf_input_r (65 downto 2)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 66;
                    when 3 =>
                        buf_input_r (66 downto 3)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 67;
                    when 4 =>
                        buf_input_r (67 downto 4)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 68;
                    when 5 =>
                        buf_input_r (68 downto 5)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 69;
                    when 6 =>
                        buf_input_r (69 downto 6)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 70;
                    when 7 =>
                        buf_input_r (70 downto 7)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 71;
                    when 8 =>
                        buf_input_r (71 downto 8)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 72;
                    when 9 =>
                        buf_input_r (72 downto 9)    <= data_in(63 downto 0);
                        bits_in_buffer               <= 73;
                    when 10 =>
                        buf_input_r (73 downto 10)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 74;
                    when 11 =>
                        buf_input_r (74 downto 11)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 75;
                    when 12 =>
                        buf_input_r (75 downto 12)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 76;
                    when 13 =>
                        buf_input_r (76 downto 13)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 77;
                    when 14 =>
                        buf_input_r (77 downto 14)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 78;
                    when 15 =>
                        buf_input_r (78 downto 15)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 79;
                    when 16 =>
                        buf_input_r (79 downto 16)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 80;
                    when 17 =>
                        buf_input_r (80 downto 17)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 81;
                    when 18 =>
                        buf_input_r (81 downto 18)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 82;
                    when 19 =>
                        buf_input_r (82 downto 19)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 83;
                    when 20 =>
                        buf_input_r (83 downto 20)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 84;
                    when 21 =>
                        buf_input_r (84 downto 21)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 85;
                    when 22 =>
                        buf_input_r (85 downto 22)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 86;
                    when 23 =>
                        buf_input_r (86 downto 23)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 87;
                    when 24 =>
                        buf_input_r (87 downto 24)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 88;
                    when 25 =>
                        buf_input_r (88 downto 25)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 89;
                    when 26 =>
                        buf_input_r (89 downto 26)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 90;
                    when 27 =>
                        buf_input_r (90 downto 27)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 91;
                    when 28 =>
                        buf_input_r (91 downto 28)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 92;
                    when 29 =>
                        buf_input_r (92 downto 29)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 93;
                    when 30 =>
                        buf_input_r (93 downto 30)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 94;
                    when 31 =>
                        buf_input_r (94 downto 31)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 95;
                    when 32 =>
                        buf_input_r (95 downto 32)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 96;
                    when 33 =>
                        buf_input_r (96 downto 33)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 97;
                    when 34 =>
                        buf_input_r (97 downto 34)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 98;
                    when 35 =>
                        buf_input_r (98 downto 35)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 99;
                    when 36 =>
                        buf_input_r (99 downto 36)   <= data_in(63 downto 0);
                        bits_in_buffer               <= 100;
                    when 37 =>
                        buf_input_r (100 downto 37)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 101;
                    when 38 =>
                        buf_input_r (101 downto 38)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 102;
                    when 39 =>
                        buf_input_r (102 downto 39)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 103;
                    when 40 =>
                        buf_input_r (103 downto 40)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 104;
                    when 41 =>
                        buf_input_r (104 downto 41)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 105;
                    when 42 =>
                        buf_input_r (105 downto 42)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 106;
                    when 43 =>
                        buf_input_r (106 downto 43)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 107;
                    when 44 =>
                        buf_input_r (107 downto 44)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 108;
                    when 45 =>
                        buf_input_r (108 downto 45)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 109;
                    when 46 =>
                        buf_input_r (109 downto 46)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 110;
                    when 47 =>
                        buf_input_r (110 downto 47)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 111;
                    when 48 =>
                        buf_input_r (111 downto 48)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 112;
                    when 49 =>
                        buf_input_r (112 downto 49)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 113;
                    when 50 =>
                        buf_input_r (113 downto 50)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 114;
                    when 51 =>
                        buf_input_r (114 downto 51)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 115;
                    when 52 =>
                        buf_input_r (115 downto 52)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 116;
                    when 53 =>
                        buf_input_r (116 downto 53)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 117;
                    when 54 =>
                        buf_input_r (117 downto 54)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 118;
                    when 55 =>
                        buf_input_r (118 downto 55)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 119;
                    when 56 =>
                        buf_input_r (119 downto 56)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 120;
                    when 57 =>
                        buf_input_r (120 downto 57)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 121;
                    when 58 =>
                        buf_input_r (121 downto 58)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 122;
                    when 59 =>
                        buf_input_r (122 downto 59)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 123;
                    when 60 =>
                        buf_input_r (123 downto 60)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 124;
                    when 61 =>
                        buf_input_r (124 downto 61)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 125;
                    when 62 =>
                        buf_input_r (125 downto 62)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 126;
                    when 63 =>
                        buf_input_r (126 downto 63)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 127;
                    when 64 =>
                        buf_input_r (127 downto 64)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 128;
                    when 65 =>
                        buf_input_r (128 downto 65)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 129;
                    when 66 =>
                        buf_input_r (129 downto 66)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 130;
                    when 67 =>
                        buf_input_r (130 downto 67)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 131;
                    when 68 =>
                        buf_input_r (131 downto 68)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 132;
                    when 69 =>
                        buf_input_r (132 downto 69)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 133;
                    when 70 =>
                        buf_input_r (133 downto 70)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 134;
                    when 71 =>
                        buf_input_r (134 downto 71)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 135;
                    when 72 =>
                        buf_input_r (135 downto 72)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 136;
                    when 73 =>
                        buf_input_r (136 downto 73)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 137;
                    when 74 =>
                        buf_input_r (137 downto 74)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 138;
                    when 75 =>
                        buf_input_r (138 downto 75)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 139;
                    when 76 =>
                        buf_input_r (139 downto 76)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 140;
                    when 77 =>
                        buf_input_r (140 downto 77)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 141;
                    when 78 =>
                        buf_input_r (141 downto 78)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 142;
                    when 79 =>
                        buf_input_r (142 downto 79)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 143;
                    when 80 =>
                        buf_input_r (143 downto 80)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 144;
                    when 81 =>
                        buf_input_r (144 downto 81)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 145;
                    when 82 =>
                        buf_input_r (145 downto 82)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 146;
                    when 83 =>
                        buf_input_r (146 downto 83)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 147;
                    when 84 =>
                        buf_input_r (147 downto 84)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 148;
                    when 85 =>
                        buf_input_r (148 downto 85)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 149;
                    when 86 =>
                        buf_input_r (149 downto 86)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 150;
                    when 87 =>
                        buf_input_r (150 downto 87)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 151;
                    when 88 =>
                        buf_input_r (151 downto 88)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 152;
                    when 89 =>
                        buf_input_r (152 downto 89)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 153;
                    when 90 =>
                        buf_input_r (153 downto 90)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 154;
                    when 91 =>
                        buf_input_r (154 downto 91)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 155;
                    when 92 =>
                        buf_input_r (155 downto 92)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 156;
                    when 93 =>
                        buf_input_r (156 downto 93)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 157;
                    when 94 =>
                        buf_input_r (157 downto 94)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 158;
                    when 95 =>
                        buf_input_r (158 downto 95)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 159;
                    when 96 =>
                        buf_input_r (159 downto 96)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 160;
                    when 97 =>
                        buf_input_r (160 downto 97)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 161;
                    when 98 =>
                        buf_input_r (161 downto 98)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 162;
                    when 99 =>
                        buf_input_r (162 downto 99)  <= data_in(63 downto 0);
                        bits_in_buffer               <= 163;
                    when 100 =>
                        buf_input_r (163 downto 100) <= data_in(63 downto 0);
                        bits_in_buffer               <= 164;
                    when 101 =>
                        buf_input_r (164 downto 101) <= data_in(63 downto 0);
                        bits_in_buffer               <= 165;
                    when 102 =>
                        buf_input_r (165 downto 102) <= data_in(63 downto 0);
                        bits_in_buffer               <= 166;
                    when 103 =>
                        buf_input_r (166 downto 103) <= data_in(63 downto 0);
                        bits_in_buffer               <= 167;
                    when 104 =>
                        buf_input_r (167 downto 104) <= data_in(63 downto 0);
                        bits_in_buffer               <= 168;
                    when 105 =>
                        buf_input_r (168 downto 105) <= data_in(63 downto 0);
                        bits_in_buffer               <= 169;
                    when 106 =>
                        buf_input_r (169 downto 106) <= data_in(63 downto 0);
                        bits_in_buffer               <= 170;
                    when 107 =>
                        buf_input_r (170 downto 107) <= data_in(63 downto 0);
                        bits_in_buffer               <= 171;
                    when 108 =>
                        buf_input_r (171 downto 108) <= data_in(63 downto 0);
                        bits_in_buffer               <= 172;
                    when 109 =>
                        buf_input_r (172 downto 109) <= data_in(63 downto 0);
                        bits_in_buffer               <= 173;
                    when 110 =>
                        buf_input_r (173 downto 110) <= data_in(63 downto 0);
                        bits_in_buffer               <= 174;
                    when 111 =>
                        buf_input_r (174 downto 111) <= data_in(63 downto 0);
                        bits_in_buffer               <= 175;
                    when 112 =>
                        buf_input_r (175 downto 112) <= data_in(63 downto 0);
                        bits_in_buffer               <= 176;
                    when 113 =>
                        buf_input_r (176 downto 113) <= data_in(63 downto 0);
                        bits_in_buffer               <= 177;
                    when 114 =>
                        buf_input_r (177 downto 114) <= data_in(63 downto 0);
                        bits_in_buffer               <= 178;
                    when 115 =>
                        buf_input_r (178 downto 115) <= data_in(63 downto 0);
                        bits_in_buffer               <= 179;
                    when 116 =>
                        buf_input_r (179 downto 116) <= data_in(63 downto 0);
                        bits_in_buffer               <= 180;
                    when 117 =>
                        buf_input_r (180 downto 117) <= data_in(63 downto 0);
                        bits_in_buffer               <= 181;
                    when 118 =>
                        buf_input_r (181 downto 118) <= data_in(63 downto 0);
                        bits_in_buffer               <= 182;
                    when 119 =>
                        buf_input_r (182 downto 119) <= data_in(63 downto 0);
                        bits_in_buffer               <= 183;
                    when 120 =>
                        buf_input_r (183 downto 120) <= data_in(63 downto 0);
                        bits_in_buffer               <= 184;
                    when 121 =>
                        buf_input_r (184 downto 121) <= data_in(63 downto 0);
                        bits_in_buffer               <= 185;
                    when 122 =>
                        buf_input_r (185 downto 122) <= data_in(63 downto 0);
                        bits_in_buffer               <= 186;
                    when 123 =>
                        buf_input_r (186 downto 123) <= data_in(63 downto 0);
                        bits_in_buffer               <= 187;
                    when 124 =>
                        buf_input_r (187 downto 124) <= data_in(63 downto 0);
                        bits_in_buffer               <= 188;
                    when 125 =>
                        buf_input_r (188 downto 125) <= data_in(63 downto 0);
                        bits_in_buffer               <= 189;
                    when 126 =>
                        buf_input_r (189 downto 126) <= data_in(63 downto 0);
                        bits_in_buffer               <= 190;
                    when 127 =>
                        buf_input_r (190 downto 127) <= data_in(63 downto 0);
                        bits_in_buffer               <= 191;
                    when 128 =>
                        buf_input_r (191 downto 128) <= data_in(63 downto 0);
                        bits_in_buffer               <= 192;
                    when 129 =>
                        buf_input_r (192 downto 129) <= data_in(63 downto 0);
                        bits_in_buffer               <= 193;
                    when 130 =>
                        buf_input_r (193 downto 130) <= data_in(63 downto 0);
                        bits_in_buffer               <= 194;
                    when 131 =>
                        buf_input_r (194 downto 131) <= data_in(63 downto 0);
                        bits_in_buffer               <= 195;
                    when 132 =>
                        buf_input_r (195 downto 132) <= data_in(63 downto 0);
                        bits_in_buffer               <= 196;
                    when 133 =>
                        buf_input_r (196 downto 133) <= data_in(63 downto 0);
                        bits_in_buffer               <= 197;
                    when 134 =>
                        buf_input_r (197 downto 134) <= data_in(63 downto 0);
                        bits_in_buffer               <= 198;
                    when 135 =>
                        buf_input_r (198 downto 135) <= data_in(63 downto 0);
                        bits_in_buffer               <= 199;
                    when 136 =>
                        buf_input_r (199 downto 136) <= data_in(63 downto 0);
                        bits_in_buffer               <= 200;
                    when 137 =>
                        buf_input_r (200 downto 137) <= data_in(63 downto 0);
                        bits_in_buffer               <= 201;
                    when 138 =>
                        buf_input_r (201 downto 138) <= data_in(63 downto 0);
                        bits_in_buffer               <= 202;
                    when 139 =>
                        buf_input_r (202 downto 139) <= data_in(63 downto 0);
                        bits_in_buffer               <= 203;
                    when 140 =>
                        buf_input_r (203 downto 140) <= data_in(63 downto 0);
                        bits_in_buffer               <= 204;
                    when 141 =>
                        buf_input_r (204 downto 141) <= data_in(63 downto 0);
                        bits_in_buffer               <= 205;
                    when 142 =>
                        buf_input_r (205 downto 142) <= data_in(63 downto 0);
                        bits_in_buffer               <= 206;
                    when 143 =>
                        buf_input_r (206 downto 143) <= data_in(63 downto 0);
                        bits_in_buffer               <= 207;
                    when 144 =>
                        buf_input_r (207 downto 144) <= data_in(63 downto 0);
                        bits_in_buffer               <= 208;
                    when 145 =>
                        buf_input_r (208 downto 145) <= data_in(63 downto 0);
                        bits_in_buffer               <= 209;
                    when 146 =>
                        buf_input_r (209 downto 146) <= data_in(63 downto 0);
                        bits_in_buffer               <= 210;
                    when 147 =>
                        buf_input_r (210 downto 147) <= data_in(63 downto 0);
                        bits_in_buffer               <= 211;
                    when 148 =>
                        buf_input_r (211 downto 148) <= data_in(63 downto 0);
                        bits_in_buffer               <= 212;
                    when 149 =>
                        buf_input_r (212 downto 149) <= data_in(63 downto 0);
                        bits_in_buffer               <= 213;
                    when 150 =>
                        buf_input_r (213 downto 150) <= data_in(63 downto 0);
                        bits_in_buffer               <= 214;
                    when 151 =>
                        buf_input_r (214 downto 151) <= data_in(63 downto 0);
                        bits_in_buffer               <= 215;
                    when 152 =>
                        buf_input_r (215 downto 152) <= data_in(63 downto 0);
                        bits_in_buffer               <= 216;
                    when 153 =>
                        buf_input_r (216 downto 153) <= data_in(63 downto 0);
                        bits_in_buffer               <= 217;
                    when 154 =>
                        buf_input_r (217 downto 154) <= data_in(63 downto 0);
                        bits_in_buffer               <= 218;
                    when 155 =>
                        buf_input_r (218 downto 155) <= data_in(63 downto 0);
                        bits_in_buffer               <= 219;
                    when 156 =>
                        buf_input_r (219 downto 156) <= data_in(63 downto 0);
                        bits_in_buffer               <= 220;
                    when 157 =>
                        buf_input_r (220 downto 157) <= data_in(63 downto 0);
                        bits_in_buffer               <= 221;
                    when 158 =>
                        buf_input_r (221 downto 158) <= data_in(63 downto 0);
                        bits_in_buffer               <= 222;
                    when 159 =>
                        buf_input_r (222 downto 159) <= data_in(63 downto 0);
                        bits_in_buffer               <= 223;
                    when 160 =>
                        buf_input_r (223 downto 160) <= data_in(63 downto 0);
                        bits_in_buffer               <= 224;
                    when 161 =>
                        buf_input_r (224 downto 161) <= data_in(63 downto 0);
                        bits_in_buffer               <= 225;
                    when 162 =>
                        buf_input_r (225 downto 162) <= data_in(63 downto 0);
                        bits_in_buffer               <= 226;
                    when 163 =>
                        buf_input_r (226 downto 163) <= data_in(63 downto 0);
                        bits_in_buffer               <= 227;
                    when 164 =>
                        buf_input_r (227 downto 164) <= data_in(63 downto 0);
                        bits_in_buffer               <= 228;
                    when 165 =>
                        buf_input_r (228 downto 165) <= data_in(63 downto 0);
                        bits_in_buffer               <= 229;
                    when 166 =>
                        buf_input_r (229 downto 166) <= data_in(63 downto 0);
                        bits_in_buffer               <= 230;
                    when 167 =>
                        buf_input_r (230 downto 167) <= data_in(63 downto 0);
                        bits_in_buffer               <= 231;
                    when 168 =>
                        buf_input_r (231 downto 168) <= data_in(63 downto 0);
                        bits_in_buffer               <= 232;
                    when 169 =>
                        buf_input_r (232 downto 169) <= data_in(63 downto 0);
                        bits_in_buffer               <= 233;
                    when 170 =>
                        buf_input_r (233 downto 170) <= data_in(63 downto 0);
                        bits_in_buffer               <= 234;
                    when 171 =>
                        buf_input_r (234 downto 171) <= data_in(63 downto 0);
                        bits_in_buffer               <= 235;
                    when 172 =>
                        buf_input_r (235 downto 172) <= data_in(63 downto 0);
                        bits_in_buffer               <= 236;
                    when 173 =>
                        buf_input_r (236 downto 173) <= data_in(63 downto 0);
                        bits_in_buffer               <= 237;
                    when 174 =>
                        buf_input_r (237 downto 174) <= data_in(63 downto 0);
                        bits_in_buffer               <= 238;
                    when 175 =>
                        buf_input_r (238 downto 175) <= data_in(63 downto 0);
                        bits_in_buffer               <= 239;
                    when 176 =>
                        buf_input_r (239 downto 176) <= data_in(63 downto 0);
                        bits_in_buffer               <= 240;
                    when 177 =>
                        buf_input_r (240 downto 177) <= data_in(63 downto 0);
                        bits_in_buffer               <= 241;
                    when 178 =>
                        buf_input_r (241 downto 178) <= data_in(63 downto 0);
                        bits_in_buffer               <= 242;
                    when 179 =>
                        buf_input_r (242 downto 179) <= data_in(63 downto 0);
                        bits_in_buffer               <= 243;
                    when 180 =>
                        buf_input_r (243 downto 180) <= data_in(63 downto 0);
                        bits_in_buffer               <= 244;
                    when 181 =>
                        buf_input_r (244 downto 181) <= data_in(63 downto 0);
                        bits_in_buffer               <= 245;
                    when 182 =>
                        buf_input_r (245 downto 182) <= data_in(63 downto 0);
                        bits_in_buffer               <= 246;
                    when 183 =>
                        buf_input_r (246 downto 183) <= data_in(63 downto 0);
                        bits_in_buffer               <= 247;
                    when 184 =>
                        buf_input_r (247 downto 184) <= data_in(63 downto 0);
                        bits_in_buffer               <= 248;
                    when 185 =>
                        buf_input_r (248 downto 185) <= data_in(63 downto 0);
                        bits_in_buffer               <= 249;
                    when 186 =>
                        buf_input_r (249 downto 186) <= data_in(63 downto 0);
                        bits_in_buffer               <= 250;
                    when 187 =>
                        buf_input_r (250 downto 187) <= data_in(63 downto 0);
                        bits_in_buffer               <= 251;
                    when 188 =>
                        buf_input_r (251 downto 188) <= data_in(63 downto 0);
                        bits_in_buffer               <= 252;
                    when 189 =>
                        buf_input_r (252 downto 189) <= data_in(63 downto 0);
                        bits_in_buffer               <= 253;
                    when 190 =>
                        buf_input_r (253 downto 190) <= data_in(63 downto 0);
                        bits_in_buffer               <= 254;
                    when 191 =>
                        buf_input_r (254 downto 191) <= data_in(63 downto 0);
                        bits_in_buffer               <= 255;
                    when 192 =>
                        buf_input_r (255 downto 192) <= data_in(63 downto 0);
                        bits_in_buffer               <= 256;
                    when 193 =>
                        buf_input_r (256 downto 193) <= data_in(63 downto 0);
                        bits_in_buffer               <= 257;
                    when 194 =>
                        buf_input_r (257 downto 194) <= data_in(63 downto 0);
                        bits_in_buffer               <= 258;
                    when 195 =>
                        buf_input_r (258 downto 195) <= data_in(63 downto 0);
                        bits_in_buffer               <= 259;
                    when 196 =>
                        buf_input_r (259 downto 196) <= data_in(63 downto 0);
                        bits_in_buffer               <= 260;
                    when 197 =>
                        buf_input_r (260 downto 197) <= data_in(63 downto 0);
                        bits_in_buffer               <= 261;
                    when 198 =>
                        buf_input_r (261 downto 198) <= data_in(63 downto 0);
                        bits_in_buffer               <= 262;
                    when 199 =>
                        buf_input_r (262 downto 199) <= data_in(63 downto 0);
                        bits_in_buffer               <= 263;
                    when 200 =>
                        buf_input_r (263 downto 200) <= data_in(63 downto 0);
                        bits_in_buffer               <= 264;
                    when 201 =>
                        buf_input_r (264 downto 201) <= data_in(63 downto 0);
                        bits_in_buffer               <= 265;
                    when 202 =>
                        buf_input_r (265 downto 202) <= data_in(63 downto 0);
                        bits_in_buffer               <= 266;
                    when 203 =>
                        buf_input_r (266 downto 203) <= data_in(63 downto 0);
                        bits_in_buffer               <= 267;
                    when 204 =>
                        buf_input_r (267 downto 204) <= data_in(63 downto 0);
                        bits_in_buffer               <= 268;
                    when 205 =>
                        buf_input_r (268 downto 205) <= data_in(63 downto 0);
                        bits_in_buffer               <= 269;
                    when 206 =>
                        buf_input_r (269 downto 206) <= data_in(63 downto 0);
                        bits_in_buffer               <= 270;
                    when 207 =>
                        buf_input_r (270 downto 207) <= data_in(63 downto 0);
                        bits_in_buffer               <= 271;
                    when 208 =>
                        buf_input_r (271 downto 208) <= data_in(63 downto 0);
                        bits_in_buffer               <= 272;
                    when 209 =>
                        buf_input_r (272 downto 209) <= data_in(63 downto 0);
                        bits_in_buffer               <= 273;
                    when 210 =>
                        buf_input_r (273 downto 210) <= data_in(63 downto 0);
                        bits_in_buffer               <= 274;
                    when 211 =>
                        buf_input_r (274 downto 211) <= data_in(63 downto 0);
                        bits_in_buffer               <= 275;
                    when 212 =>
                        buf_input_r (275 downto 212) <= data_in(63 downto 0);
                        bits_in_buffer               <= 276;
                    when 213 =>
                        buf_input_r (276 downto 213) <= data_in(63 downto 0);
                        bits_in_buffer               <= 277;
                    when 214 =>
                        buf_input_r (277 downto 214) <= data_in(63 downto 0);
                        bits_in_buffer               <= 278;
                    when 215 =>
                        buf_input_r (278 downto 215) <= data_in(63 downto 0);
                        bits_in_buffer               <= 279;
                    when 216 =>
                        buf_input_r (279 downto 216) <= data_in(63 downto 0);
                        bits_in_buffer               <= 280;
                    when 217 =>
                        buf_input_r (280 downto 217) <= data_in(63 downto 0);
                        bits_in_buffer               <= 281;
                    when 218 =>
                        buf_input_r (281 downto 218) <= data_in(63 downto 0);
                        bits_in_buffer               <= 282;
                    when 219 =>
                        buf_input_r (282 downto 219) <= data_in(63 downto 0);
                        bits_in_buffer               <= 283;
                    when 220 =>
                        buf_input_r (283 downto 220) <= data_in(63 downto 0);
                        bits_in_buffer               <= 284;
                    when 221 =>
                        buf_input_r (284 downto 221) <= data_in(63 downto 0);
                        bits_in_buffer               <= 285;
                    when 222 =>
                        buf_input_r (285 downto 222) <= data_in(63 downto 0);
                        bits_in_buffer               <= 286;
                    when 223 =>
                        buf_input_r (286 downto 223) <= data_in(63 downto 0);
                        bits_in_buffer               <= 287;
                    when 224 =>
                        buf_input_r (287 downto 224) <= data_in(63 downto 0);
                        bits_in_buffer               <= 288;
                    when 225 =>
                        buf_input_r (288 downto 225) <= data_in(63 downto 0);
                        bits_in_buffer               <= 289;
                    when 226 =>
                        buf_input_r (289 downto 226) <= data_in(63 downto 0);
                        bits_in_buffer               <= 290;
                    when 227 =>
                        buf_input_r (290 downto 227) <= data_in(63 downto 0);
                        bits_in_buffer               <= 291;
                    when 228 =>
                        buf_input_r (291 downto 228) <= data_in(63 downto 0);
                        bits_in_buffer               <= 292;
                    when 229 =>
                        buf_input_r (292 downto 229) <= data_in(63 downto 0);
                        bits_in_buffer               <= 293;
                    when 230 =>
                        buf_input_r (293 downto 230) <= data_in(63 downto 0);
                        bits_in_buffer               <= 294;
                    when 231 =>
                        buf_input_r (294 downto 231) <= data_in(63 downto 0);
                        bits_in_buffer               <= 295;
                    when 232 =>
                        buf_input_r (295 downto 232) <= data_in(63 downto 0);
                        bits_in_buffer               <= 296;
                    when 233 =>
                        buf_input_r (296 downto 233) <= data_in(63 downto 0);
                        bits_in_buffer               <= 297;
                    when 234 =>
                        buf_input_r (297 downto 234) <= data_in(63 downto 0);
                        bits_in_buffer               <= 298;
                    when 235 =>
                        buf_input_r (298 downto 235) <= data_in(63 downto 0);
                        bits_in_buffer               <= 299;
                    when 236 =>
                        buf_input_r (299 downto 236) <= data_in(63 downto 0);
                        bits_in_buffer               <= 300;
                    when 237 =>
                        buf_input_r (300 downto 237) <= data_in(63 downto 0);
                        bits_in_buffer               <= 301;
                    when 238 =>
                        buf_input_r (301 downto 238) <= data_in(63 downto 0);
                        bits_in_buffer               <= 302;
                    when 239 =>
                        buf_input_r (302 downto 239) <= data_in(63 downto 0);
                        bits_in_buffer               <= 303;
                    when 240 =>
                        buf_input_r (303 downto 240) <= data_in(63 downto 0);
                        bits_in_buffer               <= 304;
                    when 241 =>
                        buf_input_r (304 downto 241) <= data_in(63 downto 0);
                        bits_in_buffer               <= 305;
                    when 242 =>
                        buf_input_r (305 downto 242) <= data_in(63 downto 0);
                        bits_in_buffer               <= 306;
                    when 243 =>
                        buf_input_r (306 downto 243) <= data_in(63 downto 0);
                        bits_in_buffer               <= 307;
                    when 244 =>
                        buf_input_r (307 downto 244) <= data_in(63 downto 0);
                        bits_in_buffer               <= 308;
                    when 245 =>
                        buf_input_r (308 downto 245) <= data_in(63 downto 0);
                        bits_in_buffer               <= 309;
                    when 246 =>
                        buf_input_r (309 downto 246) <= data_in(63 downto 0);
                        bits_in_buffer               <= 310;
                    when 247 =>
                        buf_input_r (310 downto 247) <= data_in(63 downto 0);
                        bits_in_buffer               <= 311;
                    when 248 =>
                        buf_input_r (311 downto 248) <= data_in(63 downto 0);
                        bits_in_buffer               <= 312;
                    when 249 =>
                        buf_input_r (312 downto 249) <= data_in(63 downto 0);
                        bits_in_buffer               <= 313;
                    when 250 =>
                        buf_input_r (313 downto 250) <= data_in(63 downto 0);
                        bits_in_buffer               <= 314;
                    when 251 =>
                        buf_input_r (314 downto 251) <= data_in(63 downto 0);
                        bits_in_buffer               <= 315;
                    when 252 =>
                        buf_input_r (315 downto 252) <= data_in(63 downto 0);
                        bits_in_buffer               <= 316;
                    when 253 =>
                        buf_input_r (316 downto 253) <= data_in(63 downto 0);
                        bits_in_buffer               <= 317;
                    when 254 =>
                        buf_input_r (317 downto 254) <= data_in(63 downto 0);
                        bits_in_buffer               <= 318;
                    when 255 =>
                        buf_input_r (318 downto 255) <= data_in(63 downto 0);
                        bits_in_buffer               <= 319;
                    when 256 =>
                        buf_input_r (319 downto 256) <= data_in(63 downto 0);
                        bits_in_buffer               <= 320;
                    when 257 =>
                        buf_input_r (320 downto 257) <= data_in(63 downto 0);
                        bits_in_buffer               <= 321;
                    when 258 =>
                        buf_input_r (321 downto 258) <= data_in(63 downto 0);
                        bits_in_buffer               <= 322;
                    when 259 =>
                        buf_input_r (322 downto 259) <= data_in(63 downto 0);
                        bits_in_buffer               <= 323;
                    when 260 =>
                        buf_input_r (323 downto 260) <= data_in(63 downto 0);
                        bits_in_buffer               <= 324;
                    when 261 =>
                        buf_input_r (324 downto 261) <= data_in(63 downto 0);
                        bits_in_buffer               <= 325;
                    when 262 =>
                        buf_input_r (325 downto 262) <= data_in(63 downto 0);
                        bits_in_buffer               <= 326;
                    when 263 =>
                        buf_input_r (326 downto 263) <= data_in(63 downto 0);
                        bits_in_buffer               <= 327;
                    when 264 =>
                        buf_input_r (327 downto 264) <= data_in(63 downto 0);
                        bits_in_buffer               <= 328;
                    when 265 =>
                        buf_input_r (328 downto 265) <= data_in(63 downto 0);
                        bits_in_buffer               <= 329;
                    when 266 =>
                        buf_input_r (329 downto 266) <= data_in(63 downto 0);
                        bits_in_buffer               <= 330;
                    when 267 =>
                        buf_input_r (330 downto 267) <= data_in(63 downto 0);
                        bits_in_buffer               <= 331;
                    when 268 =>
                        buf_input_r (331 downto 268) <= data_in(63 downto 0);
                        bits_in_buffer               <= 332;
                    when 269 =>
                        buf_input_r (332 downto 269) <= data_in(63 downto 0);
                        bits_in_buffer               <= 333;
                    when 270 =>
                        buf_input_r (333 downto 270) <= data_in(63 downto 0);
                        bits_in_buffer               <= 334;
                    when 271 =>
                        buf_input_r (334 downto 271) <= data_in(63 downto 0);
                        bits_in_buffer               <= 335;
                    when 272 =>
                        buf_input_r (335 downto 272) <= data_in(63 downto 0);
                        bits_in_buffer               <= 336;
                    when 273 =>
                        buf_input_r (336 downto 273) <= data_in(63 downto 0);
                        bits_in_buffer               <= 337;
                    when 274 =>
                        buf_input_r (337 downto 274) <= data_in(63 downto 0);
                        bits_in_buffer               <= 338;
                    when 275 =>
                        buf_input_r (338 downto 275) <= data_in(63 downto 0);
                        bits_in_buffer               <= 339;
                    when 276 =>
                        buf_input_r (339 downto 276) <= data_in(63 downto 0);
                        bits_in_buffer               <= 340;
                    when 277 =>
                        buf_input_r (340 downto 277) <= data_in(63 downto 0);
                        bits_in_buffer               <= 341;
                    when 278 =>
                        buf_input_r (341 downto 278) <= data_in(63 downto 0);
                        bits_in_buffer               <= 342;
                    when 279 =>
                        buf_input_r (342 downto 279) <= data_in(63 downto 0);
                        bits_in_buffer               <= 343;
                    when 280 =>
                        buf_input_r (343 downto 280) <= data_in(63 downto 0);
                        bits_in_buffer               <= 344;
                    when 281 =>
                        buf_input_r (344 downto 281) <= data_in(63 downto 0);
                        bits_in_buffer               <= 345;
                    when 282 =>
                        buf_input_r (345 downto 282) <= data_in(63 downto 0);
                        bits_in_buffer               <= 346;
                    when 283 =>
                        buf_input_r (346 downto 283) <= data_in(63 downto 0);
                        bits_in_buffer               <= 347;
                    when 284 =>
                        buf_input_r (347 downto 284) <= data_in(63 downto 0);
                        bits_in_buffer               <= 348;
                    when 285 =>
                        buf_input_r (348 downto 285) <= data_in(63 downto 0);
                        bits_in_buffer               <= 349;
                    when 286 =>
                        buf_input_r (349 downto 286) <= data_in(63 downto 0);
                        bits_in_buffer               <= 350;
                    when 287 =>
                        buf_input_r (350 downto 287) <= data_in(63 downto 0);
                        bits_in_buffer               <= 351;
                    when 288 =>
                        buf_input_r (351 downto 288) <= data_in(63 downto 0);
                        bits_in_buffer               <= 352;
                    when 289 =>
                        buf_input_r (352 downto 289) <= data_in(63 downto 0);
                        bits_in_buffer               <= 353;
                    when 290 =>
                        buf_input_r (353 downto 290) <= data_in(63 downto 0);
                        bits_in_buffer               <= 354;
                    when 291 =>
                        buf_input_r (354 downto 291) <= data_in(63 downto 0);
                        bits_in_buffer               <= 355;
                    when 292 =>
                        buf_input_r (355 downto 292) <= data_in(63 downto 0);
                        bits_in_buffer               <= 356;
                    when 293 =>
                        buf_input_r (356 downto 293) <= data_in(63 downto 0);
                        bits_in_buffer               <= 357;
                    when 294 =>
                        buf_input_r (357 downto 294) <= data_in(63 downto 0);
                        bits_in_buffer               <= 358;
                    when 295 =>
                        buf_input_r (358 downto 295) <= data_in(63 downto 0);
                        bits_in_buffer               <= 359;
                    when 296 =>
                        buf_input_r (359 downto 296) <= data_in(63 downto 0);
                        bits_in_buffer               <= 360;
                    when 297 =>
                        buf_input_r (360 downto 297) <= data_in(63 downto 0);
                        bits_in_buffer               <= 361;
                    when 298 =>
                        buf_input_r (361 downto 298) <= data_in(63 downto 0);
                        bits_in_buffer               <= 362;
                    when 299 =>
                        buf_input_r (362 downto 299) <= data_in(63 downto 0);
                        bits_in_buffer               <= 363;
                    when 300 =>
                        buf_input_r (363 downto 300) <= data_in(63 downto 0);
                        bits_in_buffer               <= 364;
                    when 301 =>
                        buf_input_r (364 downto 301) <= data_in(63 downto 0);
                        bits_in_buffer               <= 365;
                    when 302 =>
                        buf_input_r (365 downto 302) <= data_in(63 downto 0);
                        bits_in_buffer               <= 366;
                    when 303 =>
                        buf_input_r (366 downto 303) <= data_in(63 downto 0);
                        bits_in_buffer               <= 367;
                    when 304 =>
                        buf_input_r (367 downto 304) <= data_in(63 downto 0);
                        bits_in_buffer               <= 368;
                    when 305 =>
                        buf_input_r (368 downto 305) <= data_in(63 downto 0);
                        bits_in_buffer               <= 369;
                    when 306 =>
                        buf_input_r (369 downto 306) <= data_in(63 downto 0);
                        bits_in_buffer               <= 370;
                    when 307 =>
                        buf_input_r (370 downto 307) <= data_in(63 downto 0);
                        bits_in_buffer               <= 371;
                    when 308 =>
                        buf_input_r (371 downto 308) <= data_in(63 downto 0);
                        bits_in_buffer               <= 372;
                    when 309 =>
                        buf_input_r (372 downto 309) <= data_in(63 downto 0);
                        bits_in_buffer               <= 373;
                    when 310 =>
                        buf_input_r (373 downto 310) <= data_in(63 downto 0);
                        bits_in_buffer               <= 374;
                    when 311 =>
                        buf_input_r (374 downto 311) <= data_in(63 downto 0);
                        bits_in_buffer               <= 375;
                    when 312 =>
                        buf_input_r (375 downto 312) <= data_in(63 downto 0);
                        bits_in_buffer               <= 376;
                    when 313 =>
                        buf_input_r (376 downto 313) <= data_in(63 downto 0);
                        bits_in_buffer               <= 377;
                    when 314 =>
                        buf_input_r (377 downto 314) <= data_in(63 downto 0);
                        bits_in_buffer               <= 378;
                    when 315 =>
                        buf_input_r (378 downto 315) <= data_in(63 downto 0);
                        bits_in_buffer               <= 379;
                    when 316 =>
                        buf_input_r (379 downto 316) <= data_in(63 downto 0);
                        bits_in_buffer               <= 380;
                    when 317 =>
                        buf_input_r (380 downto 317) <= data_in(63 downto 0);
                        bits_in_buffer               <= 381;
                    when 318 =>
                        buf_input_r (381 downto 318) <= data_in(63 downto 0);
                        bits_in_buffer               <= 382;
                    when 319 =>
                        buf_input_r (382 downto 319) <= data_in(63 downto 0);
                        bits_in_buffer               <= 383;
                    when 320 =>
                        buf_input_r (383 downto 320) <= data_in(63 downto 0);
                        bits_in_buffer               <= 384;
                    when 321 =>
                        buf_input_r (384 downto 321) <= data_in(63 downto 0);
                        bits_in_buffer               <= 385;
                    when 322 =>
                        buf_input_r (385 downto 322) <= data_in(63 downto 0);
                        bits_in_buffer               <= 386;
                    when 323 =>
                        buf_input_r (386 downto 323) <= data_in(63 downto 0);
                        bits_in_buffer               <= 387;
                    when 324 =>
                        buf_input_r (387 downto 324) <= data_in(63 downto 0);
                        bits_in_buffer               <= 388;
                    when 325 =>
                        buf_input_r (388 downto 325) <= data_in(63 downto 0);
                        bits_in_buffer               <= 389;
                    when 326 =>
                        buf_input_r (389 downto 326) <= data_in(63 downto 0);
                        bits_in_buffer               <= 390;
                    when 327 =>
                        buf_input_r (390 downto 327) <= data_in(63 downto 0);
                        bits_in_buffer               <= 391;
                    when 328 =>
                        buf_input_r (391 downto 328) <= data_in(63 downto 0);
                        bits_in_buffer               <= 392;
                    when 329 =>
                        buf_input_r (392 downto 329) <= data_in(63 downto 0);
                        bits_in_buffer               <= 393;
                    when 330 =>
                        buf_input_r (393 downto 330) <= data_in(63 downto 0);
                        bits_in_buffer               <= 394;
                    when 331 =>
                        buf_input_r (394 downto 331) <= data_in(63 downto 0);
                        bits_in_buffer               <= 395;
                    when 332 =>
                        buf_input_r (395 downto 332) <= data_in(63 downto 0);
                        bits_in_buffer               <= 396;
                    when 333 =>
                        buf_input_r (396 downto 333) <= data_in(63 downto 0);
                        bits_in_buffer               <= 397;
                    when 334 =>
                        buf_input_r (397 downto 334) <= data_in(63 downto 0);
                        bits_in_buffer               <= 398;
                    when 335 =>
                        buf_input_r (398 downto 335) <= data_in(63 downto 0);
                        bits_in_buffer               <= 399;
                    when 336 =>
                        buf_input_r (399 downto 336) <= data_in(63 downto 0);
                        bits_in_buffer               <= 400;
                    when 337 =>
                        buf_input_r (400 downto 337) <= data_in(63 downto 0);
                        bits_in_buffer               <= 401;
                    when 338 =>
                        buf_input_r (401 downto 338) <= data_in(63 downto 0);
                        bits_in_buffer               <= 402;
                    when 339 =>
                        buf_input_r (402 downto 339) <= data_in(63 downto 0);
                        bits_in_buffer               <= 403;
                    when 340 =>
                        buf_input_r (403 downto 340) <= data_in(63 downto 0);
                        bits_in_buffer               <= 404;
                    when 341 =>
                        buf_input_r (404 downto 341) <= data_in(63 downto 0);
                        bits_in_buffer               <= 405;
                    when 342 =>
                        buf_input_r (405 downto 342) <= data_in(63 downto 0);
                        bits_in_buffer               <= 406;
                    when 343 =>
                        buf_input_r (406 downto 343) <= data_in(63 downto 0);
                        bits_in_buffer               <= 407;
                    when 344 =>
                        buf_input_r (407 downto 344) <= data_in(63 downto 0);
                        bits_in_buffer               <= 408;
                    when 345 =>
                        buf_input_r (408 downto 345) <= data_in(63 downto 0);
                        bits_in_buffer               <= 409;
                    when 346 =>
                        buf_input_r (409 downto 346) <= data_in(63 downto 0);
                        bits_in_buffer               <= 410;
                    when 347 =>
                        buf_input_r (410 downto 347) <= data_in(63 downto 0);
                        bits_in_buffer               <= 411;
                    when 348 =>
                        buf_input_r (411 downto 348) <= data_in(63 downto 0);
                        bits_in_buffer               <= 412;
                    when 349 =>
                        buf_input_r (412 downto 349) <= data_in(63 downto 0);
                        bits_in_buffer               <= 413;
                    when 350 =>
                        buf_input_r (413 downto 350) <= data_in(63 downto 0);
                        bits_in_buffer               <= 414;
                    when 351 =>
                        buf_input_r (414 downto 351) <= data_in(63 downto 0);
                        bits_in_buffer               <= 415;
                    when 352 =>
                        buf_input_r (415 downto 352) <= data_in(63 downto 0);
                        bits_in_buffer               <= 416;
                    when 353 =>
                        buf_input_r (416 downto 353) <= data_in(63 downto 0);
                        bits_in_buffer               <= 417;
                    when 354 =>
                        buf_input_r (417 downto 354) <= data_in(63 downto 0);
                        bits_in_buffer               <= 418;
                    when 355 =>
                        buf_input_r (418 downto 355) <= data_in(63 downto 0);
                        bits_in_buffer               <= 419;
                    when 356 =>
                        buf_input_r (419 downto 356) <= data_in(63 downto 0);
                        bits_in_buffer               <= 420;
                    when 357 =>
                        buf_input_r (420 downto 357) <= data_in(63 downto 0);
                        bits_in_buffer               <= 421;
                    when 358 =>
                        buf_input_r (421 downto 358) <= data_in(63 downto 0);
                        bits_in_buffer               <= 422;
                    when 359 =>
                        buf_input_r (422 downto 359) <= data_in(63 downto 0);
                        bits_in_buffer               <= 423;
                    when 360 =>
                        buf_input_r (423 downto 360) <= data_in(63 downto 0);
                        bits_in_buffer               <= 424;
                    when 361 =>
                        buf_input_r (424 downto 361) <= data_in(63 downto 0);
                        bits_in_buffer               <= 425;
                    when 362 =>
                        buf_input_r (425 downto 362) <= data_in(63 downto 0);
                        bits_in_buffer               <= 426;
                    when 363 =>
                        buf_input_r (426 downto 363) <= data_in(63 downto 0);
                        bits_in_buffer               <= 427;
                    when 364 =>
                        buf_input_r (427 downto 364) <= data_in(63 downto 0);
                        bits_in_buffer               <= 428;
                    when 365 =>
                        buf_input_r (428 downto 365) <= data_in(63 downto 0);
                        bits_in_buffer               <= 429;
                    when 366 =>
                        buf_input_r (429 downto 366) <= data_in(63 downto 0);
                        bits_in_buffer               <= 430;
                    when 367 =>
                        buf_input_r (430 downto 367) <= data_in(63 downto 0);
                        bits_in_buffer               <= 431;
                    when 368 =>
                        buf_input_r (431 downto 368) <= data_in(63 downto 0);
                        bits_in_buffer               <= 432;
                    when 369 =>
                        buf_input_r (432 downto 369) <= data_in(63 downto 0);
                        bits_in_buffer               <= 433;
                    when 370 =>
                        buf_input_r (433 downto 370) <= data_in(63 downto 0);
                        bits_in_buffer               <= 434;
                    when 371 =>
                        buf_input_r (434 downto 371) <= data_in(63 downto 0);
                        bits_in_buffer               <= 435;
                    when 372 =>
                        buf_input_r (435 downto 372) <= data_in(63 downto 0);
                        bits_in_buffer               <= 436;
                    when 373 =>
                        buf_input_r (436 downto 373) <= data_in(63 downto 0);
                        bits_in_buffer               <= 437;
                    when 374 =>
                        buf_input_r (437 downto 374) <= data_in(63 downto 0);
                        bits_in_buffer               <= 438;
                    when 375 =>
                        buf_input_r (438 downto 375) <= data_in(63 downto 0);
                        bits_in_buffer               <= 439;
                    when 376 =>
                        buf_input_r (439 downto 376) <= data_in(63 downto 0);
                        bits_in_buffer               <= 440;
                    when 377 =>
                        buf_input_r (440 downto 377) <= data_in(63 downto 0);
                        bits_in_buffer               <= 441;
                    when 378 =>
                        buf_input_r (441 downto 378) <= data_in(63 downto 0);
                        bits_in_buffer               <= 442;
                    when 379 =>
                        buf_input_r (442 downto 379) <= data_in(63 downto 0);
                        bits_in_buffer               <= 443;
                    when 380 =>
                        buf_input_r (443 downto 380) <= data_in(63 downto 0);
                        bits_in_buffer               <= 444;
                    when 381 =>
                        buf_input_r (444 downto 381) <= data_in(63 downto 0);
                        bits_in_buffer               <= 445;
                    when 382 =>
                        buf_input_r (445 downto 382) <= data_in(63 downto 0);
                        bits_in_buffer               <= 446;
                    when 383 =>
                        buf_input_r (446 downto 383) <= data_in(63 downto 0);
                        bits_in_buffer               <= 447;
                    when 384 =>
                        buf_input_r (447 downto 384) <= data_in(63 downto 0);
                        bits_in_buffer               <= 448;
                    when 385 =>
                        buf_input_r (448 downto 385) <= data_in(63 downto 0);
                        bits_in_buffer               <= 449;
                    when 386 =>
                        buf_input_r (449 downto 386) <= data_in(63 downto 0);
                        bits_in_buffer               <= 450;
                    when 387 =>
                        buf_input_r (450 downto 387) <= data_in(63 downto 0);
                        bits_in_buffer               <= 451;
                    when 388 =>
                        buf_input_r (451 downto 388) <= data_in(63 downto 0);
                        bits_in_buffer               <= 452;
                    when 389 =>
                        buf_input_r (452 downto 389) <= data_in(63 downto 0);
                        bits_in_buffer               <= 453;
                    when 390 =>
                        buf_input_r (453 downto 390) <= data_in(63 downto 0);
                        bits_in_buffer               <= 454;
                    when 391 =>
                        buf_input_r (454 downto 391) <= data_in(63 downto 0);
                        bits_in_buffer               <= 455;
                    when 392 =>
                        buf_input_r (455 downto 392) <= data_in(63 downto 0);
                        bits_in_buffer               <= 456;
                    when 393 =>
                        buf_input_r (456 downto 393) <= data_in(63 downto 0);
                        bits_in_buffer               <= 457;
                    when 394 =>
                        buf_input_r (457 downto 394) <= data_in(63 downto 0);
                        bits_in_buffer               <= 458;
                    when 395 =>
                        buf_input_r (458 downto 395) <= data_in(63 downto 0);
                        bits_in_buffer               <= 459;
                    when 396 =>
                        buf_input_r (459 downto 396) <= data_in(63 downto 0);
                        bits_in_buffer               <= 460;
                    when 397 =>
                        buf_input_r (460 downto 397) <= data_in(63 downto 0);
                        bits_in_buffer               <= 461;
                    when 398 =>
                        buf_input_r (461 downto 398) <= data_in(63 downto 0);
                        bits_in_buffer               <= 462;
                    when 399 =>
                        buf_input_r (462 downto 399) <= data_in(63 downto 0);
                        bits_in_buffer               <= 463;
                    when 400 =>
                        buf_input_r (463 downto 400) <= data_in(63 downto 0);
                        bits_in_buffer               <= 464;
                    when 401 =>
                        buf_input_r (464 downto 401) <= data_in(63 downto 0);
                        bits_in_buffer               <= 465;
                    when 402 =>
                        buf_input_r (465 downto 402) <= data_in(63 downto 0);
                        bits_in_buffer               <= 466;
                    when 403 =>
                        buf_input_r (466 downto 403) <= data_in(63 downto 0);
                        bits_in_buffer               <= 467;
                    when 404 =>
                        buf_input_r (467 downto 404) <= data_in(63 downto 0);
                        bits_in_buffer               <= 468;
                    when 405 =>
                        buf_input_r (468 downto 405) <= data_in(63 downto 0);
                        bits_in_buffer               <= 469;
                    when 406 =>
                        buf_input_r (469 downto 406) <= data_in(63 downto 0);
                        bits_in_buffer               <= 470;
                    when 407 =>
                        buf_input_r (470 downto 407) <= data_in(63 downto 0);
                        bits_in_buffer               <= 471;
                    when 408 =>
                        buf_input_r (471 downto 408) <= data_in(63 downto 0);
                        bits_in_buffer               <= 472;
                    when 409 =>
                        buf_input_r (472 downto 409) <= data_in(63 downto 0);
                        bits_in_buffer               <= 473;
                    when 410 =>
                        buf_input_r (473 downto 410) <= data_in(63 downto 0);
                        bits_in_buffer               <= 474;
                    when 411 =>
                        buf_input_r (474 downto 411) <= data_in(63 downto 0);
                        bits_in_buffer               <= 475;
                    when 412 =>
                        buf_input_r (475 downto 412) <= data_in(63 downto 0);
                        bits_in_buffer               <= 476;
                    when 413 =>
                        buf_input_r (476 downto 413) <= data_in(63 downto 0);
                        bits_in_buffer               <= 477;
                    when 414 =>
                        buf_input_r (477 downto 414) <= data_in(63 downto 0);
                        bits_in_buffer               <= 478;
                    when 415 =>
                        buf_input_r (478 downto 415) <= data_in(63 downto 0);
                        bits_in_buffer               <= 479;
                    when 416 =>
                        buf_input_r (479 downto 416) <= data_in(63 downto 0);
                        bits_in_buffer               <= 480;
                    when 417 =>
                        buf_input_r (480 downto 417) <= data_in(63 downto 0);
                        bits_in_buffer               <= 481;
                    when 418 =>
                        buf_input_r (481 downto 418) <= data_in(63 downto 0);
                        bits_in_buffer               <= 482;
                    when 419 =>
                        buf_input_r (482 downto 419) <= data_in(63 downto 0);
                        bits_in_buffer               <= 483;
                    when 420 =>
                        buf_input_r (483 downto 420) <= data_in(63 downto 0);
                        bits_in_buffer               <= 484;
                    when 421 =>
                        buf_input_r (484 downto 421) <= data_in(63 downto 0);
                        bits_in_buffer               <= 485;
                    when 422 =>
                        buf_input_r (485 downto 422) <= data_in(63 downto 0);
                        bits_in_buffer               <= 486;
                    when 423 =>
                        buf_input_r (486 downto 423) <= data_in(63 downto 0);
                        bits_in_buffer               <= 487;
                    when 424 =>
                        buf_input_r (487 downto 424) <= data_in(63 downto 0);
                        bits_in_buffer               <= 488;
                    when 425 =>
                        buf_input_r (488 downto 425) <= data_in(63 downto 0);
                        bits_in_buffer               <= 489;
                    when 426 =>
                        buf_input_r (489 downto 426) <= data_in(63 downto 0);
                        bits_in_buffer               <= 490;
                    when 427 =>
                        buf_input_r (490 downto 427) <= data_in(63 downto 0);
                        bits_in_buffer               <= 491;
                    when 428 =>
                        buf_input_r (491 downto 428) <= data_in(63 downto 0);
                        bits_in_buffer               <= 492;
                    when others =>
                end case;
            end if;
        --else
                --out_rdy_r <= '0';
        end if;
    end if;
end process;
end arch_word_expander_64IN_to_493OUT;